��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O���kâUP	~NS��O�Irb�c��\<��⺧A
��Lr��'&ageY��7y�4�}H�&ˊt������[	Ni?��^P��R8Q�P0�B͍Y��y:�eDM'��}�r�S�N���m����>��af:�@����3�݂���V�I�z6�0���EI]��0Z,kPD#��u1��!1>`=���3�e�#��|��.^(�Tmh�|��k�����t֦,�V��� ]U���
2i찻���ڇҚ�����"(7CyK�ox�Da�:�7�V��[��I� �hy��n]{�v�kV���F5K�q��~*���w@(:ص�O_Ok�g����R�~�g���5�i5�sT� ^xL0�1�oR���HŅC���u�鹰��TЇ>A\!�fP/���Gt��5l�r3��FՆc?jR�R�N��k�R���_��G3�؟��B"ei�c�CT��"�D��8��zwIne��]�0-S��"����a��Y@����*Q�Nu���:_�/]3����HT
�$���"�	{In� �=<�Y��٨}��M����M-�:gO�|��rS����H`�%����ᵜj�%��|P�d_��r��wwc�06�`V�	UA��h���$6@
����� ~�l��b���z�����l�U�6��Y��7����-�y��L'U��yb���{��(pW����3����O����ˑ��� �ʻ)A���V�#���)�q |g|�M̙UQ��H�vB�
��q������=|~P�C��!���u?�9e��