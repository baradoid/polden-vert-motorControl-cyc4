��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�=l��!ӻ���C�&�m���bݧ�5���iL^�o��ȿ�T�*rʇ���q�-G~�&S�P�	�A��J����b;��QUU�;�%��R�Ǻ�(�	��F���CŔ����!�,d���+��5JZ���F�q>�6�xp���,���\q�l���4�"4�d|�kn�F�B
1qv�T�ۉAD��iQ$d���ĸ�餋6t� ��byE诫G����}���o�S�T-*f��loo��M|M��攛䑼4��:F��<����ɇ���%��O��/�׸�3����E�� �.�-�E
���h}�3a-�s)m�^��gKJ����d��)�Xus+�a�̺ej��2�b>5�D���1��h/�U�m>0��w{Ӄ}������u?���h`��1�)�5� �huDo�Q�-�N�M'"Eb��CzfA.V�j�b=I$Є֦���n�5O�ǫ`�==��x�8$y���䇛h��_��67����k�#�}�z�9k �&��u7
c�2��K'�/�xq�c�{?v\ą���k^1gG3{�}K�0�A2���.� �1g�Y��IfͩF�Pt���ظE�3�J^���j��d��%_��x-?A#f*>7�����uW�V����\�u��4G�w���5��W��{��A�n[�l����p�4ͬR,C�~J �B^�5Y�v^��W��I��rbV�h����cr��1��B��(�n׵��q/%b��=l�j�bg Q��z��<���NoBx�y]Y�&6�l8<��f�N���O��_��	)Yԩ^Ɋ*��4hx�٘|�~k�.�HN�E "uu�!�MFr%���Xq����(+�1Pw� S��T�:��:3���J@f#0�U��'�W�>��'2����
����I<J�Ь~�ǰG�i��/�ɘ�x��OJ��ID�������%�!���F�����]+�g��je!� �L��<�`E����]�'e������+Nr��������Q0%Qh�3�.h�X�lom�{sn�6D�L<�+1�f��=�K�x�۝�rЕ�%�w8~���G�Eg��ǫ �O�6����!%� ���b��o*�up?�a�W���䚯y��@�$��!R�*�e�)KYG,�,�