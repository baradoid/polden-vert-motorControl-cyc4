��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��[���G�8��2��}>���=��Ó��>�	�E�fr�p̮=�@�hӠ�s\\p[ �}S|�.������M��~��c�\�Pf���0x:aV��{�5Hk
��V;F>O\U���c��ML��!�XcNU�fXR;^R��tn$�c�#�}�H�&�3�)�txG`)���Cv�->|��(��J��6:_�{��,��x���(/��4@������NW���x�܎�Ȳۼ`������Qz�sX�zjtB#Etu���M�0�h�g�*���ֱ��@q��׳��l�C }���j���!�0
̚d�l�""a�lՄ 8�?������n\�;��IiP�@r,��ja6Xa�4L��^�Ԧ���&k�q0�	9S�	F
;��M��ܚ�=��@�����r?�-���$����y@_Їo���~4��:�YB��v�l#�"�cO�/�ә{��-�e�K��?�X��P^#R$<���,�ܜO������i��"V��}ȥL�ɐy2W�rr��^���7��yu^�>�5)ۋ,���>b��,%m���,yS{�^�_k�mAl���0�̃ԩ�+%��h�J񶩗텏���|�J���p0e��E��J�z���r��,lIp1"9GՋ���ҹ&\	"���N��,4�O��PJ��j������]0�	����w�M1�������-#�
t0$�_���\�w8�ہ�t���{�'���9�W}7z��6�����ڰ|T� 2'��D �zb��V�\�g@��Ki��5	�c��$S�r��oRctLBV�!�Iᯆ)�ilc��5Ѭ��p���sj��7p�G��T�*�d8������qM��� Z�������_�c��,i�(92dWE���Zzo�2�6b���{s�eۅeK�맅T��Q��I�µS��Tuw�؊	�֗��
����?�T�~擨b.���Ҁ�`3��T�4MJ�J�����?w�ItZQG��K��灛SH`�S�����8�=h��~[=��x��
NB��gɈ�yt�(�P�p�� &�dn,`�D���R<k>�c7U��o����;
:�tԑ&x���n��?!��KX��T%K�m����u��������Nc�ʢ��9NUD ~��N`�͎��Ѩ�����$�+��
pOç�\��c�B��Cy1��Jq�w���f���tI�>~�oV��s�^��5>�� �i�"���9hJ��r��u �!~niE7f�V�E�1O�F;x��]�e .�n4� �:�sЍǭ��/���\���>#����e6惩l'P�yz�z���N��ّ�����;C�2�Q.R��By͍�	���^E@�j��H�a�%�[l�o�q�,��mU(�`��o����y"*u57�Ni�/�Wd�~�ۙ[��)�AV�M��GJ9c�VD��7�7�ph�������XՊ�pky�C�>�(\�Ri��&�WG�U��^�k��ר˓[�����T'�m���)4]�~"l-�p��/_�@�V��p�oO�����1�fզY5�^������wCxbL�R�B���9�i?�G��^i$����Bf�w�ԛ+�7ρI��=���aג�C����g��%5����ލ�J`�'|Ds�PD����A��x�	�P�B� Ð�n�����E�dK|KZz�#R�4���\���}���ʗu&'��!�ھYO�� !���-~���6+`Q54���ҕ�~��@�����
��p옻0uT;D���(<��T�\s�3睙 �Y�ba,-���1� �Z�,�ܼ�D��1#������z�tON?C�h>�~o������O4I/�I�qe�7qQ����;����d��ˬ����;�dVcM��]Unv;ߋ���u#;߆<g̔1tr�.����<�D�(ɓ�T.�����w�#�N�TQ��I�k��Y���@v3���5�8Ҍ���=O�"ĤJ]�(T2�go�,��t�U�9����ʹ)K֒���i��f���
����D�g��H��VJ	���Bg9yb ���q*�-?��b"<��C�����خ<�LvRO�tk�C�(C�t���O N�g�"/�3/��,/~=���
�q>�ޚ���apN��	ǅc������>6m��Q��\k1�+'&8�*!���Ov+!頉Z���g��"�ﺍ'�k&�Vy�q���1��M��3<2����Lh����\�ty6m�[LFV�Ɓ����ߺ�b4�nF���������}bΌK���n�t�C�w#I�s�VQ�~�M>Vh���j���L��,[��uF+k$g���Z�Bf�[~�p�yDFie�]l'����Y��;�D���t٫W�{��$`�O��?P��:�Zϋ��x�i���A�D�$�n>��j��~��֔f�b,n�`�h9
��c �M�@0w|��ƚ}3k�����/�Y��u�i����d�2���L r�6�;\�+�_᳉��x�`��OFY�Y���!���������/�p���?]��d;�=��}�o�2d�{�P�>3e^�j�kq�P�(4�Uc�Dڵ!:�Տ��T�ۛ��n�~I��.	�����Xrۓ�3eI&5��MVn	����<Co�>RH�sr��%�ev�m��рu�š�������o*�D�^�iU\{ċ`	LF�0-0^dV���H����I?�� i�`r�j����Hv�w�䁙s��`J=^���+�y�2Տ�vg`c�����W#��L�.���LF-�,�j �K�����xB����A�@x��ʘ��'* t�z���F�	����'����"�X3%|�SA�X{R���{�g0��	�9u��P�q�w��P�e�ERmH��Sz�Ww�ۣ�
��?j1� ��v�i�('�+hd��r=0�c�alr�a�~m[�q+��B��r��d�簎���<}��ӄ?%m)'ڍw�YqxrO�Jd�]P�о��<�E���hP�T���I0�HSZŌB+���#@�~��0�ni�#Ǉ�n0���=�29ޭMUX�'����@�|ϧ5�܁�L1S͊��G�iL������G���_b'Ƭ�a h���4��kʏ� l<@���a�7����W��z�(�l�+Ο�&�C����?}\�ک�?�}���v�ٿ�)	��#�іi���N)��!5���%c��dk`W�A��^���.6_����!����\5P)'Tb3��F����?��}��k�����C)G�Y���'+0��n�1����fE�!�c&�6s�}���W�<�>Z�"�iSa���_|��0۷�k=�k����b?shYZ�e9[��ؒ�A��dd������tz��a���l�~,�`�',��޸/�V���/:�̫%_y��
����?�Tྮ��G��\�;g��k�sC�0�]��Lӕ�����K���������1k��ʊn헙t)������8�6���:���q���*�ky�s�Ю, O_���]��r����G�G�ʘ�jYb+��c���	���8�4zhqCf}	Q1��_aw�0�,F�� X�#�DJ:�ϒP����Wl��'����9��8$��:<KT�Cq�������&���Q�L���<�t�"q��������%�ݜ����ܸo�����R�����*a���G��^�b�����y�}�J+�u�:{M �T��<0Te!��O˷�.y�wnner�����@���=���G>��4g1�7.�?�u��F�VV���A�k�	�-J���NZsH��	Amľ��>�c��� 9K�@�T�E�ׂb�����:	���pxSn�+YYx:^YR䭶�ؖ��,"��R�bՎ���h��թ��Y�����G�j�M/@\&��SJ���NÁ�K�9�>f%�a�9Ǜ"�Ȋ$M9�)3����sYc�c+֢�OYN��Nm\��86u�n�	%�3�~n�?�"�����0�R`�/'d`��"�q�l��K�`���