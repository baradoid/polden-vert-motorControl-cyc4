��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�H]�0��L���V��&ZF��C��o<�2��ߣ׳��J7������B��2�%�Z�����dњ��P=f�uq1�cdcэ��եѵ��y|Ty,�*0�ߊV���FRA�p
/98k��Y�U�5SR����#""�'��up��;�2��aO�i �0"X5�;#�g}м�aX18� �,���NgB���nN�EK�qӋt�1�/c���I�N�L���x
�0�_�CO�
�z�F�v3R��`_:@񜾤5�ѳ
�׫G�5АuPH�b)��mH�^ehV�/�	$�X*��\.�;򿜵�p���+�ހ��2� &�ʿ')��z�E��'I|�0"��׶��L�b��-[���=���<�MO0ʗj�k�WoQ �S��Ҿ?d�Hs�[Xf#�N|�K�⑕�e�N�ݘ�҈���ڲͥ=�U,*��Ҋ������}���\q< 3���k�,T��8��8+Ă��dG5��4	����j)?��գ��RV�GIb�4�e �.;��4C�EF�J,g��Ĩ����y��pUӈ?��֧�[g)�;<�wK��
�Y>�kJ�f�Q vO�7�*��L��H��C/�H�[� e��V���}��N�2ML�u�fyt�N�W���G�T�����%z����6�e@�����v7�?l���wœ���0i���mNtoN�
�F{��kڗ�LH�|`�k;����~�]�0-�������������e@�=�p���)\I��Wi�a��O�����_�5J㤠���w�T�VV�g%��6����xn���\':י�n�B���H�1:F�\���3RM��O{��	�*�}#C��"�7�"ָ<)�tn�NB [<���L;�h\x�!s�Ⱦ���gE�;���ܩ!:|��"!�l|�gm��=D�@��,�Cxi�j�3�o�]/<��1R�?��|�?[����ks����St:���Q�L�}����?��ܶ�����Ә��;��ã����H�� k��#������~8`�)�@���6��e�Rw� P&x�$����� �ٻ�u_wt�K�O��+L`xe�S����o�*����|��}q��3ũ�,��U�Q�G	��=VUZ���7d�ܔx� ��|A�s���G�����C]�r�� U���Mhz�ұ�F��z��"��EAU��rJvx ���!VeX1���k@1!��5�6��	�2���yMa����y�_�G���4�V`�I�P����MZ*Q.к�ĳg�Z�������������
�%]��{��;Dx�N?��p���*�Y��2��,_��o�������ݒ�\pq��U����˷�W6<��۝�,��~s��$�"ᩬ�g����t��t�F� �N����&�\�^�+$kw��pq-Ӏ�&'J�K2�݂�>�h��-�|`��N���3��,� �̈́�jYV4S��:��s��'��L�)��9P�J(��87�s ���Z�v
<��|�L�ߪ�z-�>�D|ZI��2���9��Uh����"�6��3��r����"W��@�o�{�~�hT�?�e�U���]�O�d7Vi��c���K�L �Y�u����\&I���Dmd&�&���{,��X������K�o�z�1ؒ��߁�����?'Ċ��ڻȌ��8�FE�S���} l�\���d�h�Kw�y0F�.����0���X��I�*�J����B��g19��CW c�_�wepr*3�r�@�z����s,'c�j�FZ��4�ȟ��������{�ʻ(٬����X;?�iϮ$IN�s �R�
���>��a���us5�c������C�7�{�������^Bh��}��;\���&WKG����U�@��57�l��DK�pX�{��2(���G:�d����=���Ap�!P�#���n�zŔ�>��,D��{Sv@�)�R11	4Q	��u?�\��1��v���&qlH�p�>sT�	�I^�9vmՁ��6Q���|��n.a�OTh�!V��?�	��K��Wܶ[;)S�:��d��rt=v��RE��_W���Q����*x�o������ʬ�{���z��A;��� �W�Wt ��]�U���2K��孯$;?~�@�X�g��"��W+;+"$Si��I5�C�Y���Z�,V�����6��@Y�xk�>.��#���n��j
s/PT�;߶��}��)l�Ĉ���ˀ�!���[�v郚�J����bR.��9h�l��\�]�&�ވ�@�'W����;v����BɶIg@�Y��q��[�T���D���n�x�#[��h\���0��m�g"K���<�im;�(���6Uט�0.���":ھ`-�
�!�����]��Bw�M�2��ۥ�#VW������iI�� ���X �Z�_�C�o�V!ę�����kЗ��V��]֕��cv��6��M�L���p1�`��K�J��L1ɠ�y�#��l�(�$� �c��������~CG�������OM@��6��ƅ<�,E��4aؖf��W.ˢ"��Gj<�P����(��D�ǣ�	 (����q�>���^lU�D��C���J���Y*����l�x������a�>��)��9έC6��	S�C���-:��X��C�7��x�<�_�Ӫq7	�s���i�y� -%�f�X��t+�w��>L�]�����ԛu�`zQŠ�P���`��OJ���_'RxZ췑"x�ywX�Ҥ��㍕uA��*�u������D�%МLy��H{p���4(��c �$x�p҃����HI�������^&A�
��쫋{٤�j�W� ���di�1[�x��l�?N���7��}�@m����>�C���쵏�ޘ�L�<$D��a��C����2�k�Q�sQ�\�͑��\-V��1kv�d��ɜv�nw�u��V���Y�`�nO.�k1�Υ�V?E������=���Β��#��������