��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�
#��.{и�5��+d�N�~�>ve��Pp��$���n�_g	�%��y�a���ۋ%�E?⻁�T���P{�3��9�)=�� ýDd^ǽ����
��N0��g�횅::R�[(W�Y�o�js͎pĎ�҇��w1�l�e7��P��)�]�Z[���|����������m*س˥�q�j���t�Lq���.@����ۦf�}I21����o��ۮDmT�A�ģ~��۷�|��)�(z+����g�M(����.�hZ9ؤ�%��C��df����UU8�C9e���rH��5)�ט�F����OV	�r�8��e@T���c[����~b*��<P3�\�i1ڦD6����PX��>}�l�_[�j���؞!��/������r�%]e�s�[:mH���q��W0Ʀu�@���Ԑ�AU
b��4@eE��Re^r�������r_���vi�83E�:p�R�/2��B��Iw��u2$�=�-�Գ�6.�wI^�#WN� ��� �4��u�Z$~J�� �[2T	~D���=����u@s��4_�����bv��7%؅��K���"c�KqxW�W�d��!1й�����Ő!�0S
c��[���\���Ķ�l�2N���+��� 3ۋ�����,�[D_��	���dO�qX����l��Hأ4�Y �}.B���2s��g�����F;��f�j�!Z���p�e+�MR;������H��W��� _�t\�nB4��`�02u��t��
�ϲ��o s ڤ��01�Q	��x��?�uH �87�szj�B�à�Z��1d�p�q����b~�z����Y����Z|$��&���˚����� ��XK�I� i೟�[�ʋRZ�N�u&��H��.?��f�A9�1Q�>�8�}�Cߛ����iQ'L�:۠0�7��$ǩd��2Qi�5�rOZ��5��c!�����IG1
�O�i��4����M��Bx$�B���F���S��_|��	�r�R�G1񘀝<���L��П����CV���h�BjC]5��|�^K��. ˓_3�K�]8
c�>�-��Q��&��̈����Ud#���݃DF��/�2x/1Q�h�#��<.#���:~Z�S���l����-){�Lj�G�[���C*�D��t!«����i��������l )+j��&l�)D��y�"s[�	� 2x-l�|Z��"?'r�5��^���!��6�A��e��	�{�Q_l�k�f�<�:ɷ�����������R�]:
/2v˽m蕉�	�i�3`ϑ���b͙d�0�v�8(�T*�h�i�]��f��"���/Q0�>V4箑.�@�V9i�Z�c�1i�A'~nz�˜����I����͛�=�M��h.F���n .[:���E���M�vq?���k��T_k��b�*�+uL�Ԧ|������(n�+y7��WǸ������fFO"� d�o)�p����76��}�)���޶4���ӽS������K�s�W�\�0M�ʔez�Ɛ�N��{�^G�)��LI�~S'������k3gt�~�������@)]��h����2���Juע��X���&P�c���,c`�ѳe'����~V��ZL�yG?���!i�x�zN�j{��Kʕ�P�+1���|��iȔd��<<���:s�^8E�Df��+�S-X!�a  |c��r��5+ͷ���SY�݊\+w+�/��,�u��B�� Ę�@k�	X�0�כ�?�K�N���ޮ��oыI����
BK|sslWf]��ǍavxIsx��`��ۇ���wL����O)�m=��|�*M�����0|)-���^C	�M�i��wSDff�`�T����Ԉ�\H�TU ��a�Y��� h|>?�u`���
�p�p�<��+2�i�!J���������j�-]E.�_1�?^��+�`�+��ABE��Ex �q����*%��㱮�AݱK�VDDB�]�3d��P Ow	*�՚it��m��6"Yt�ǥ�bI{� r{���Qct9��<����̰|,�!8���2����t�K��9��aaMt?�q��W<�d�Z��)'|KH���I �$����ח7z�@���.e�����_�5?|ck�
1���+�x��Q1c�8�̾Ȳ�;�׽7>d����-f��=��f�j>�����`	=9]')�.[���ϓ;��)L�EB��A������/SY�{\�`��R�P���]��uv��H
�׮�a�lZC�]������M-S�3u}�J�}�h��U�OT�ҵm;��%�/Q�q;&���d�[�y�)_�7]��^���`�����!x�`2��Y���3�ءz����C��� c�uʄ#3��Nx�z�*������b�?6#���ĂT�[`���<	P���E��˿�2N9�n��ӾXp�[��r[�)��wX����h7ȿ~�.Q�]����iq�Y��`�e8iEhp�j���K1ܺ�<u�/��U��~���'rWR���18�e�w�8�֝,���8�[�5�C����ɻ
�t��Cز'�t�-�u�A1֬�6� ���JB=��ˬl��Y-~��9C�]��2�Ӭڌ�{�.f���&gˎ�1�$p\fS���o�h�4 �Z��`"\�c�^E?�$��c ��(n�B�<}b��e��꜔e�/����UҢ�%�����׎o7��0_(�=v-U�ٓ#'�p��	�
�d5d��V�2Ơ�e�8��>Ի>�l��o#�RQK��Ʉs RB��D��'�KFn&b�e-��EiO��"R���oY�Vc�Y���C��ʳSt�cXm����za|6dĥ�M�#x��i���U�z�[])��r�(7A�]\ˈ���C!�\Q\��hX�Ah��J�i��
���KZ��E� /��gn0z�"~�no��Ia>	f4��L�,�Y�k���I\��R��B�l�����Ȗq-����q� � �cl%�ǑV�폙��imS���ߵLMb/���)ٜxs��OH���]zme��_KfFd���j8H�IM=�B���1��a��tJ1$.gu۶T� �r���5�w4�U�n6&!��G��6���J"�R�g����j��rd*�6�W���[��cm�;>{"TxC2%*N���43h��wh��܃��lo�