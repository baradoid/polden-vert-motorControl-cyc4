��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�
#��.{и��k��x��ZB�E�a���Ҕi�G4���h�#�~H�:I.��D=�0�}H��|F�b�j;���D:G��1�=0�s<�I�Db�.��,�H����i�j���t��G�G!>�����祗a�t�o�c	�zn�(e����A���(~qjׇnH	D��!�r��rn0��A*S1��1ѫƖ%�n$6e�NAֲ�;��u���������@��Y^e���J�a�:��qɎ��OJ��=�_(:A���%�wL��|�{ƚ��&0��5��`��"'�{�����̽��d>q��.�IA=g��::���R��X������S��&9e�ْ�t�|�x5�͙����b|nQL�	�Le���#�f-�7H�ּ�^�����o�2:g�E��=%�9�k/��h�*J"�k�7\fR���/~F���)�@�]�y�y�'�e��Q���ׁ�9۽��ZA�իs	��`��%�?�m�ہ�؏�<���n'/�+s̠�5	/X�EhٕG�#_��NW�:�|�����k�{�tQi��)��fzE��Ft5~_��jY��c�{�k^[hkm,`k&͜"-.j[����5Ő�G���q����BG6	K���j��e� �Q����o_K!�$�\.=X0n��>�l� �@����$�W�[$R��Uӌ�Nq�\�����"~e���5���)5� �PN_�(��T�<�~���W�26���C%1aȨ Z�f(�q\�k1��e�X�dZ�yM���$���>F��1f���I`D�xv�6�3���PM��;�	2G�id�L�����`����- ؏�L�:�LJEs'��W�'Q�T��n���m�ana9Q��۝����%�J���Jz���{5��Ӏ���+؃�����.O���s�.�#��Ӕ�yk�)Y���a-�s���-$JF����t��TM��D^c�l�R/�ҝ� =?_ʄgT��|���eZW��cY����i3h�g�
b��e���R�3O�&�]���Ѐ��'5ɩ`ޯ�Q�A��r��^���F�Sn�a�za߸�Þ.A)�KqD*���i'����pn=��>4�֤Ă(�2�8�a���]�F��� Ii�Cw}ol�����`���>�O�����̂�V�U,�L*��!�qeB�^Do����qP�]��a�ApFgߥ�k� �+�HhP�W�� �^�oF-��.l',8Fq���iW 
�L��*_�r0�G�� 5���A��X9�l��8	��+R+{S�M���qR��vq�$�l�G�ZWn��4�l�A)��w�c��^M�e�*gעҔ�U�`�s�L|���M��蘁����;~)a���dV���/�a	��� n�^����	��c8�Z�xRX�$� O��U�8w�"Լ2u>EN�b3�~�F�O�����յ���§p,R��(gY|p�C!���]bE�\�u�d��.-�a~�kL�7f�RD����m�����SHjVʦ�~O����I���j��i=��/�=0>�S���:��RH��=�K;��y����˞���G/�,��#�4CZ3ѿThE �|��
������B|��X�#�T�!��u��9j��?"u�`"�K�B�����r�׉�vm1���5|{]#i,O�ʦwf-�-�m����iG��Yg����he�O}�taA:8�(*N�楦XMG������eiačx�`pҝZ���hA�Ca&=B"+�ީ{gxm2���,It3�tqUԉX��;����  ��P�"3©�]
T�N�؈���f�ˠ�+G�ÛEa��T=� ��Z<c%���Z<8�w�k��)�n὞%��[+q�l��K���)	���7�G�t�n��I��z���4F"_8OPek���K�4�3^�\X�eA��e��:U+�!��<��j��ݣ�.����a��8tV"��@A��(��������K~mqRe+ֳd� �yO.��d.��#z���������TqEBA�Ň����������!By���𢙧t�&����fE��_��%�{���}-�	�]���<�+F�NK�|�Uk�i`d���^�)��w<�����s�hŠ*�ͫ��,6��2t~�M�Q��{�B��>ꪣDYע��G�\ip���6�N��z�f�`FM߮w�6��7�F=��H��f��\�S檷�Dع���_Ȁ��B��遈�%��9��ߴUu!Qf�B�/�
;X�C�j�̓���v���9k(��^�V�s������f3�z]��&o��s�H�~��W2�w�MN�������y�b�֒�k='q�4�H��!Q�-5��|�U�8P��r�Wy��'ہ;m���S��3��A�_D�.zEc���q�iU*LS�7���(�s?|�ZuԎ�	�D|{��+��:n�T���@M0å�̙]r�;iq���M��DɎ�Ϭ�]�s�zN�|<�)���M
O��a�۝��"{i��I��~u�ux��ͦ9�*������\��;��u�R��u�g���q�Ǚe���JbGt(g+��}����ӄ���O�{������)�'t|V���"w2�@o�����n>�z].�;�,��T��$�J��1����{�T�a~9�ˆ���G=h���r��7��6J9cb�Ph>�7�P�p��͕,�k�S�h�'�	�טp�iԏsz8��7Sq,E f�=�:�G�{&#[ΨE�ba�N})+G�+�F�{�a)�m$��jm*� �ԆP���s�mP�7�����+��E�f{�"�
���Q��V�L�R�yЂ�[qX�p�gU��+�i�{7hg��o6�!��{F����ALQ�-���q�9�c\9�pTm��Q�"o����v��\�l�w�\o�W͚��mJ9X/Ϥ+�ۮ���_��	�Ч%���+�����3�V�wT��v��C�c���/�o0d�7��m���bɠU#bz(V%W��LDq�-��Yb�Hƽ���-��#�N/�� F/˻��\�����uS$d�Ր��L�|�]�-F���ObB�m�g�����$y�I�z�UU�R���IN)wF���Vb4�t��jf� ��υ���'���k�0T���C�� G������>��N�]����ql��ز��1�uGdq��z9�մp�Qf#���3hoP�J��-�� ����F�S���nb|�pJ�A�ڻb\�tc	ɢHHTrq�	Z9bq>��� ���gb��CԥN�r骋�<���`�YO8�ji�)M�۝5�D�F�O^@2������VL\R�	�W%yޣ������h��t}�%��@D��f�*By�٨+�;O]-v���	r�j���f5���]Y�ޫa��R�EW��u|����K�&����Ra��
o$'�$?�uo8��\=�{L�x�2uA�	y�]�u��5���A����7���1�gK�)�+�Le3Ix-���3��`GP����mƛ|A�zҷv����	�9�\ܱ��,�������q;����=�U7lf�深��P|�L��6'��s '��am&9��GkTY�1wIR�4K�;~�j}ά0�~�����S3���0�|��Y��j�"�C8r#+o��2A�36���ʴM�K>7q#l�N�[������$b���6���� !�	z��bP��?a��K����y�Z�