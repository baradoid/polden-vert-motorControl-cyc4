��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�h�d�'��Ƚo�f8V��Gt'1A�S#��� ��O�'.�v�F�F�`D���:(��$x�gQ�U�T�ù)Vhs�s.�����)��L����-!������J	�E:�-�����t.V\D"�BARG�4�e^��4����ZUC�DS1_�E���i.4��_h��#n�t���"��Mtb���p�$m�_����� l�� Z�@Ur&��t՟�e5�?{��l�o<'��Y�1�PfMn	���S�����R�d���_Hz��D�#�������c����"���`�;q��M�|��O��DV�Fؿ�h��X|#��{v�
ߓ;�G7�4��L�l ��aV\Y�"�J��ڶ�Ց�
�y��z�I�t���('��v���u~rSg���`V��cih�vǄ 1�͊��	����X�)�f�K��2�w#Z�(�nj���{E'c�J9'_O6�zCa>5��;��t���=��b#(����,�L���4���B�FƩ.��7֊�y��vN�$�O�n��3eV�V�@
�2\�~��[7(�`:�	��/W
�5�;Xcy�s��x���H�����n#�D�5;���Q�JR�X����e8-Z@�T��I<k��JN
0��~=�K��>~���]��)g;X��t5v��7��+ӿ~.Ρ�kW��t; �G�{v?��J�P҃�bΡ/e ��<Ã�v���ZqC,��a����T�^�7*���u�w���A��G�cxvar�ʚ���ɖI��*ۚ}O��a敵ɛ!Ɠ��ԤT#�i��7B'O[Z񥮩z�� V�D�H�>���YX�����+��T?�7agy\*Y���� X.^�+�����U�H����	 �[�0v�Z "�\���KN\�)�"�Z4���W��I,�aK�Ұۆ���2��g2�I���p��X�����