��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�rܹ�U����<Z���mZ���hM,Ҋ����� hv��7��0��o�'p��5Q6ՙTo��cAO?8��t��1�ZH�?��"S��w�����uʻv>	8:�6���x��c�A��S]Ƨ�Bt���!�1�*֋� �smC�L�L�����F�R���`���#���|�S�&`'m��OXHu�.*��я�+(�Y��<#�Ht����ف8K�{k?�7yI�E��r�S[eK����u�lVW�o&�a\�YG���^�m���ݞHß-��R�����O#,f)ZH"ymTb��/~��j�S�.Ό#�'�j|��6��C?�S��3y$�����U�,���]�G��؇O;׫�+�K�ĕ��*Ky�00k/��ch�!��H �AcA�F�l��{T���(ٽ�vD�h';KAHz��W0ř�M���AsxC��9��̥#�ϔ|^�>xLd��LZ��A�Ӑ�Ke�[�{�	t��>OD���B�Ì�K��q"(�6�������	����Z9 ������U�;c7}p��M=[�֛��kE.@P%-���ї�J�7�$�IWT'�Z�@�	��>���p��l='⅖(}����K��ʢf �Տ����g�fcj�Nd�#��jn�C��U룲�J�<Ls�������BlP?�Dg��*��@�(�?���� �x��[��ـj�b`�pdt���`�����)/(��K�Q�S���z��R���H����2�<�zC.���5P�N�<�MY-�W8�#�H���ƍv��D�@�ɵ�-��$&R�<�{�AI��U�>J70l�W���m��J+7���-�$���Tܘz>P6 1Bq�s�~&9�d��7u�����@�����Y�$Kϓ���PH��V���>X�?�Nڢ�̤�qL۸��ެu���*�(-�#hW�Lt�� B�����>����z�>H�
.�>��Uq��HI�\s`[���Lm��5���>�\�uo�ޗe�$C�]�RO4-l
���.��{���b;�j\��t�d�69��>�@��iH�Y�J#>�hB)E�tN���3�|o ��]�ᵺr�Of�́�!���^�U�/ͥ��i�T�
���O�Rϵ��V���dS���N��(�mY$���&�Qvُ��Enl��ёΫ�T���Y[��/m�UƳ