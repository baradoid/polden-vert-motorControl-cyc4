��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�
#��.{и�9�o�FԤC�!�6-</�`I�'�U���V�B�pk�$G��|N��h�$W�n�8��}(�dO���p�+������e���A���SQ�6V'biW��$�!�~X�x��0�x�W�-�02�xO�[Į
��ϵW���I}z�*��,���G>& ���'1��@�~6&�Y!�?�8g�D(\��wn2�JV��Oy]� -��6]>ER)jr5��"���.�vߐ�|\0c]E�#�|B�B���sVЋp��G�A�n?���b���:���-��m��0��F��>��!~f������)YO#F`Zz䮙G�d]j�_!�V��pv�����VWD�,)�Ye~g�EKU �L)~�Wgp��?�S�m(y9(�Q?7}g�d��
�t�[��/Q�W�Q�`�F8eL޿���ss�-�6�Mo��+4���Ӗ��rPg-���g�~cO��yX��t;�U��p�?RL�.�
��%2����+
���}%�7��C����f�]��:��a���ڵZ)J��e$w��������d�F
�)��N�i�K��am(�ڃ�n�����E�'��	p&(��*99�4��
=��.�TΔ��zp�CK�Y��E4z�r��"k���z�C��P� `�n9�c���#-� ���Gra]��g���pd�ɟ�e�8��׺�˞�A���w��WA��N����l�[�v�3q�
�noT;k��(�|}��bM�v���:	��̴�Nt���yq��5��W����L���"3���J�юbl+:jWA�h�)c��m�o��4�6z����Ch]h�lR��Z,�ӎ�PE���_�8�v�O��a�J(��a*RG��o�w�Z�e%۹�\��A�����S�Xr�5,�].`�g�|ȫbW��� *���c�����g�	c�KzD$i�|����[�Y#�-��"�&��_K�'�\����n�0~��ՁtGrh�P��P�FQ�F�oR��v�E���A���J�V�>i��^�*�lR!S�x�\��z�b@��$��������L�:�6���`2V���C�a�$��f��rˍ���yn�32רr��F��>x�O}]��: wB��rV��nɣ�=a|}*�'|^��d��*�tPfϙ�^J��N��C���b~���86�e�ξ�2���t	A���8�d�բ�-��N��|oi��Pqk��MdȂW��6ZyQ?t��I0Aw��먝C�N|�1��`���1�6@Η�����?�n"W��C����9��tś�F��a���#�M���U�#Pw�]���c�+�ҁ�ĉl��2=�����g=��%4Ѻ_��7�-���
�'J?g6}7����h]�_j�C���_��ı��P2
:�?|�s2�i�rc���Z�_�/��C���,��\e��6���o��SF�|��ٍ����U8T�H�>��X��}s6S�[+���õ%l'yY�P�����qb�����q}�2�M��n|��E�'א��A3p�b�D��`j��-�؞ǣ����|3�;��F�C�@)o��	��>|��/gXCL�����Cсe�#9�z��@ �Bgn�x]pWT���p��V/��%t���KTCM���H�&�C$�	Ƌ>��,���e+�V��I/�1�>0!�c��ɏ.���ٓ%l��L��b��85om\@suAB�L���*�~}�?c�M�	�H[=����B�fko�����*���JD�~�L40|]oe���g��;�#F.l���y�=������A������U��'����:��;:�����Xm��;��~ϡD��%_��(��/�2Y�A�;�~t��T���ܢ�Q���I[Q��.���z�����n����I�^��%�k�k�Y�Gx>�_;��`)`��ea]� ���e���,��mK(dp'_�����4�F���CGphPy;�+�_B��^VgU�>6�K@}�H�.L����h�<b�yB���k?~�m��xkOd��8n���O�LM�-%��5��,g���LZ��C��b֏�..Z�.�H�y>Xt����灤��Q�a��1� �Itf ���Ģ���3�Tـ��-�ɱ����vd���OQ1Q��aӼ�NJ��N"D��'�X�P��K<��fHf���������v�j���*`h>�k�b'�:���Mȵ���X�0�>�b�P���HS�.@�mK-�����N9��Z���$虷ck����hq$|y�l�*l�"�1ry15�=h�m�\�
(KA��vM��t\y%'��i�B�3$�z��X�9���Nׁi��_�V*��:��5+i3��X���{$�o��Q,�>�t���ZJg!�Cΰ�,�j�{��d���?�����eͿ;1z�Xn�j��u��%�N2a�C���Lf����"���\�|�3�u�)�Z���9C9{Z�%�N�P��j/����a��"3�xL�=��ycA�O������[�̰�y�}���P�N�Ie�����#���K ���W�O��˴jit�Y����?)8�t��N؊�}E���v\B7�3��;�J�`>������`��ae��ە=l8��'w��F+���_��n��x\�T�w�CC���^��vR���a��j��t�I�����P��ma1�R��f�����rd����P�3~q��e@H91Ǿ�?;Rd�8��K�j�j�ں�����c)��rKU�����L��
S�g�2m�3��2�Q��qn�߅> #���6�� ���u��E���EA���E"EM�AC�j��˂���~���"[3D��i:��s��*����G���=Z�P>fSk2Șt�	�@;��G�mQ���N�%t!R����5�P�tχI��'� tV�qI�(��}�.+f��Ǭ�}��Q��ԭ��*��:���9�i��w��������	�d�E[���_�����<V���4J0��30�_�̥T�~�쿀�K�W�'2�H���@��D_�Ԓ��9:�Wz� b��}C�+���N�����>����At��3��7���6�J����j\gkr5�%�,��a��`��i4��$�S�����d����Q�A�k��K���Q�{����������䡳!��/�!�j�.���].ֈ��*��+�@��ߑ��p�ax-��x��=(kA&҃��_D'E�3ٜ�E�y���M<Ձ됭���B�-��O�| �:��8$��I��C��K�X1�Σ�`�PJ^~ʻ���)�R�D?wx�䮃��;c��l��pG¾�fB��e�,����	/�쓾�\�:����l��}j��n�e,nr����C��Il+k�,w��"��`)F�h]X⒨X��c�"�s����E�5K��ְo+W��}�:
���DD�%f��<G�Z�	�������O��T�a;/�+eKs����;'F�o�)�m�&M:m�"�p.ױ��l�롲accB�Ù�q�߆��/��L/�z�u?�`L"7�e�s1���F�ݏlq�P�* %+iC��0Y
�aA�@G�L	%mq���]/��uЌ\�&�\���J�}�����I����5o�s���O��d��mo�8J�̤�Wí�aʞ���Hݨ�f&���6����d�A�l/��}�>�ʹβ��%
�kБ�����g�z��7�BU�px4�R-�����`N׺�&�[�Ɏ­X.'fpE�����C�.x��D����_�#��gv�.��q��j]��n�+����':��1kPlh���d_b%���ULNB����j��#N�x#o���
�U�m��j�kqPz�/-Z���і�<�Ts7	�͢%Q?'¸}�9p�j�L�s�c�/����~��9#��`��A'-��wR�4�����~����|���[�J<Nx�|6�.s|.�{��Kf#���.Tf��VVO������
��R�c6RԕͿ̣��{R��tP�~B� ��ȝb��/�zy����3e􁓡E!;� �".���+���Ȁ�5��@�0h߭��
K��Q@� =�
�Y�틌O֙��K�)4�?IT#�dН.��������C͊;k����.�C ��H�-���0J�z@�K�!wNI���s���}Z��q�5&��"�<�S8�0�$��8����Łht����z�g�bDP[#��s��/k��X�]ΐ��[n%�<�nnH��Z]ށ���6�C��D䐮�?�@y{a�_/�}(]������7����>J�4"����o��I���Q��v�܌�[�%�v9���e��ؤ4����Jk�0o����7�
f�e���D�?��\Ntp.3(���F�p��S���k��qmX�g��m¢�u��F�*��<����葋F�Z'p:IL�?���hP}����k�&1 �䒂����b�$ҹ@��7� ë�l��\SS�������f��@ҹ0�K$g���b��cR�#J�i��3�qEqy�t��:��%.Đ�����Ì$�9؃#�AN����^��>
�\6bP��]/�X ���Ӛ���1fb[�)(��B�:��Ԉi�����%�;Tmy�Z��\f�$�]�F�g,!�.#]O�gS$w���I!��r�$� �$�3�|�_���qB>�xr��b��@�q���k)�>%�t0wPSl�?���_ 0���!uOA�dMC(w�rx5;�� �h�,����'v�G={TE�32��;Û���f;byT&eƯ�ڐ��N���:��_NcI��������7�������9