��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O���kâU���c'O)UG��t}�K�_��s�V�.��3�����xB��<��8�
�z�%$|(�������R��tfև {�U�>Ƃ�py�}X�c���5�x�`������`���5�J�@�h��ց��9.�/��ڷ��R|�u˘���3�?r����T�P�q5���w�2 ��g1~�t��)(�J�3:���$�h�V�Rm�dh���M�Sl��6�#�����T��0��:��N.��i.�����d"�.������b	�K�i(j{ܨ.��-�Q�ʇ�
9JG�*�
E�g�%���u$�m�P�L&z�)���{��LI���Ëu�Lu�7C���0�g;a��\�',ё��q��E�!�XZ��':�1���W��p%@=��~:�a�1ND��ސ���Oڶty��ɡ�HB<]BQ�8�J�-8�^fv�C�'Y��'�s�ˡ��A�����c���>=�)�@J26*�GuB��JiA�����H���|
��j�uU
.�,���(P@ޠcD��R(�d�.ڱ����L������CΥAX"�ࣽ{�:v_�/���I7���[DOy�C~%�����5���+���i�j?.i#�U~�R�6u�[��}+�qK�F���=X:��x��s�u�
GE�ѫ-� fm�����
���5	����Y鋧<�[(i�8��i��[�*��)�hCm*�=�f��|�u6���$�F,����-7a\ճb#%��o��k}>�D��
��9��;�y�육`e'D��<t�!�H�6�*�(�{ɄD���&�d| ��g�#Q���͍$"9�K�ꚲMN�T������'aoX"j�\I��Ev�s��Y�@���Ǯ(��NF7n��j���������{S����������d�'�+5�s�}N� $��꠫Zp4�iF ���AH�����U���!�:��!���@�Au�:����V���_+�z��/{ڃ����_�H�=�)"���ҧ#si'��<^��a[�IK،���e»�i�w��ުͅ4\��;S��,E�mױ%��d�W�j��9k���_zc�%i�������Ex#l�o� �M���x����)��>+w-'�������E;3: $IB��c�� �Ϡ�\x�m�q�.@������Keߤ%�ԥv*�p��C@�W5�bC�.�Ev��᡻vr�WP����:=��WC����~2A��n�;(�/�m�I-���8 �1������>��]���.����e~�iWS��9���h�2�!#\��a9�����󥨌xE���F�L��Ʃ[i"O Y&1Z걒�BW�IS��$�e�&쁜1%���9����(Ehi�{ӏ��M�3J	]����T�k������cG9)5��Q���0e�D�×�'�[<��;�S4}��W�yL���ȯ����B��.���^�DZ���>��̛��}&���!����Kᅴ���k�rm��|ӎ���QG��G��N=�]�;t�.�wT�W��lW<:DP�@=�LRcV��vd����u���T�R���)8Kh���l�Y��0UM�(�=�,�
$�
��5�_�S����2c�Ig��Q��L�%m
C#�$kn�����ۂ;�836�*3�!�����a�k��Y�o��\�:ۺ��p񃭲��j��!�fVTXc���Q8�`�6��۶3F�Z1�!F3 ���Q0�S w���%�&��o�M6���'Mcxf���
���Rb�
71������J�~���Z����C�ɏ5��Tmꋳ�YvQT;0���l��ީ�����P �`نG���KG#�1[��A���:�z[}�W;H ~��X�>e���O�h�Fس@`�B��~+/Ym�� ��p#d+)2���"c�.� ���je�$��"����Qif�g\��U�h1|��J���
���+~*���k��\��ޚG]�n�?�h�n�������^4�c���?h���`%ݦe�x�?Z�o�0�"c!3Ŷ�3~�~�ki�� 	H���1'i �]AXJG�`�Eђ�Y�CLm�C" L')���]��+,B��X\����T�z�D�G�T�^��YD���6P��}��f �C���eU Ӑ��q |f~R��Ht*g
��Z��i�|�tJ:��p4����-r
�
��eC����2�_[��uBQ�2��*H�]n��u���?m�@GD�t��3p霠 �^=S��,��E���x2�ؗ�6u?�='��a��Z��4�%�5T�e��k�x���%��[J�W\�j��@k���b���qb���{�B+�K�r7e +�'����J7����`jD����k��	S���Z�:��a�����xU&]+���`��R.!�����f�}��������_;��,&,�}��u\�*�,��%2�w��:m'BnZ���@�;�9�����n�X)�����j7Tz�k�3�GӔ�b���@�o<�|2�yzЮO�v�@���k��H��;�"fT*���<�j����A%��O+��Q�:	�^>,
k��]��j�=m�1�o�r�R�ʇt����de� �dj����F��N���{��x3��6)���fb�-4a]X��S�${ص=�A_2�zi�v����<�4�C�/o�����<��v�KHz��~��EZ�R�0K`� �j4l��|��0i�`I�������|Z�U`���j�
py��	eS2���e# pT�	on����`�l�9�b8�5�)s|�7�`��Ȣ�o�K�:����.q���;<�����y�CD��K�F���`7�>x+a�c:ܵ~�QQ���U��h}O~E��
 %v��m����:DC�#���'Z�R�`���z�=�ħ"��6O#: �~c�̊���/%�S��@	r�ʮˇ������J�o�[:�����cP�q���η��7��p���褖Ր��y��*�Ht-x!�����`�M�2�g54")��yIeȻCy��4MT%�������9����лkOOZ�]�n�\�^Z~^��2�L��ݟɁ7�=��F䖤��X�[΀��Ć�Oqhc��X�r�?�G'�Ru�N���¾�=3��+��gxhc8k�*���y3/Q�ט�3���o�!�,[�P��n#/��{m+HR��7>"���J�R>�#nI���l�C�t��G陸9�2=�O��O���tSG �AI� &��K�(���6T�d\8m�}9�Շ�T���;˯�]%����*�p�P�`�De.���4�z�9�];X:�w2�Z����f�ˡ���x:���K֚s����oF2�0B��|��}��|P��J�ՠ��4��Me�?