��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�
#��.{и�5��+d�f�&�ʬ�N�>ȉ-�A�⊓4�n,*V��'Ӿ���(����И�g�h��7�U�WYg��-���U�b�^���#���z��6�����5=LX<�6���������-�n?Q�YȜXRQ}�b��f"��h(���g��b��y���䇅�Of��}�J�&��ƌ �<�;�yn��;���c�E?�]�٬eE���q;O���|��02H�aGN~;ݥ���icSóD���<�fx�;��V-׾+����W:;!݀�A��x5�mKke�Co��V��cut�&9�W�ȡ��i�Hր��8m38�/U-5p�j��+@�a�����dW�
�<#�����W�)r(L6������Gj���aM��cK>�����;��)��m���xZ
�uC����'vA,?��(��E�ɴ�{Ԅ���<E�\�n�e
���z���]�1�f8���.̅	P������s �9grA�Y� �B�%Q@���տBT�l�r����#<A��^���LE��P}�N�L�8-Sp��Ft�!��8��f�W��Fڍ$�P����ң}����5P�D�����')��ŗ��������F@��tY"��B��w�F��d��@g^��µǃPW��aN'ť���k��~[)���  ���E�m���Yk2^&�a��qK�6h��	6a,Ts��H`�-��xA���$.ͷ��&�I��gׂ1������z���+���P�%A�,�F<|A��E�[���B�x'�?�̵�������Ā�_BD�����Tq!�|1��FO瓌�z�V`�Gx��Tj�jf}W�QI�������B�e9�Ѧ�b�* A��@j�5i��+
8��40�`-3_�����wq�m�Ͷ+���ҿ},Gv2�gC�Gs���B81)�ŧ�����z!�bc|G�A�^%l�ɪ)t����_�
>�/$�6�i¼? ����h�mI�q�S�k[�:"�5O)���Q{����`1V?Ǥ1g=��B��TU!�~�9�軐���[�)�dU䑍YOP ��Q�8ȗe��Is�;
	��(���}BM8㥘вG���j�]T;�c5Eu�E+�>Ă�ˬ�(B'�P!|��gen�Q�����UHa�7����p�A@��0��J�(��-*��毯�(I�<��g�� ��z6;� &��Ğ�OD���D�+\�袷�N�wI�U��<z�έyX���?u�l�ɒ����p�%��$4u@����퇞�)�wk�I��<�����l6�Z�3�(��DC��ޘ�+4~���-�Q��U5������&b��B�׃}&0���T��M�17SiqhrN<ZR%R3T���z��	qÇ��뾑�r�/v�{$�̝�Tr�B��r�ǟa/8h<>G�	��z�l NZ�׾������C
�8���eRt[J���V�<gySE��Y��l�~��l� ����7�sl챤4�ܬ���HN�^
�d� �x�g���;������@��m걹��4GUvع�[�a�����I�Ԗ�W�ηP�� ,�N��yX�r��VR�'X�ww�Ӑs�v-^;�X8��{Gt��.'�0z��y��ڠ&jur�[���:z0Y��A�Zb71���%�������J�l�=6�h��ّi��SS���B�&(�=�7:�vvQ��Td�Q����9�9O�#4]IH��z`O
������� 2Cn�O����J��sx�N�a�ڧ��d�"����"p}����\�{�ȓ$[�sF�I{�|�3���' �6��Ќg�͠�I���������Gٲh
S3�R�%�3a��_�!�-<v٦��gLB>]�Y�>�m�U�hY���J��2��)�G49.bxX��,�5���B������٪FG`�vXs��p��MǼ8��wy�w��E�ef�]ߥz�?��i�о�$�p��u��~�;�J�R�"�7׻��!�2粁v��K�#�-�ɉ�:0�휮��.TP�N��۬KY�?��N�.�Y���,��)��T��KR\�1-������3�\��s?M�:	2x��3��a ϵ�O8 ߊ~LT�&K;��5VЇ*���;_��v\�;��?Ў�iE�������AF'�:"|ߧ�k����>,�����,V��8Y<m�;�Fg�<H�I�+b%���ex�*��_�{�ԴSk�1�!N���Z��~z���-*?8 ��!Y�[�m�?�{��� ME�b�4wV�k9���@Kt�KחS���I��L�!Xp�ig�v%��(I�g��oM�F��V���y<X�)i0{~��A~����S�7��7��cf���[2T����gK�d�"���%�f2{/��A(b�_$���O�(ܱ��-�i�P�o�'�[4����~�W�jF�==ߑ�6&���q$