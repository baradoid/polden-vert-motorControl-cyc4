��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��[���2���W�G����-������Y�R�jZ�O�H�ȗ}�ІKʵ*�"�d���-�l�3l�%$B�F9�V/�:��`#a}TQ���A�wf�E.n�B<�l�p�g;D@������!�):dAY�zd=�N� `6d	B�zSXve\Z֋@��>���USm�u	��@�'��!2�a��U�����a�����1U�>Xbp�1Jx%{6�7�FV��{/���H�.�l>d��_���i�f���Q�g�T����M��'��"8P.�L��Ir��z����ϣV�.�L�Lo�oX���F�\�FdI#߬g��u�Osv�������( )] �B�]H���F��i�c:٩��;�0���j/���O�R����'SiA�4t�A���JNO����xj�ۿ�(����:���k�1���k ���^��6���ٿ��c��@���\�s.,�*��d��<;ټ�k�|��h���>J�D�W�k��矔҅�:��3�0ץ]k�����֣:'j��ģ'��-�)7}�9�r(J�Z�)�&���g�9D!�
7rm,�:� s�=�ho���7�(��9�l�5�פԥ��ms��iJ�	z�ҁ���@)b��c�%�/ŉ� H�!t3�`��^�a��\`3V�OgS+�@�PP��	�["A���4I��˼I�0�k����oКK�81�s�u��Ycz��e�� Ϲqv>��hKa�	w�k��Qr����)J��܎�����8'L�ܲB�1�a�v�{,9u�:1����z��꾝tI�A�֋��+Ǜ�����ZJ&ԃV�r'#W2���j�xD��C�c|kߌhF�n�9��y��?�Z�y��h�p��b��
xh�]��w�k��+9AႆA��9��B��99�gy&�
�z K���H�zd;���.�n���(31��3�4��?tco�x�f��0(����W��H/x��̀K~a���je8�/���Q����R��� �.R�KvFƻ����ʠ5b�V�,+�t)}�D|�iT��z�St�4�O��NAӸ�Y��hqSQ0NwP��y���UʳT8Qu�G/iR�:�N�R�)]��(*�"l�o��6 t���U��Ƞ^� k]����F2;��F.~r_��[��M��%?i��jy��[`�<>���%�z|���Y['-�o~@�t�Xۯ���R�����q�
.�5��A\:�;�6��3�o6��<f8C[�H��[��B��!о���P���0Ǐ��:C+���^���f��?Ɔ^��x��e7`��HM@ŤW�tA��W�d��D ��q�F��<w�uK�fW _c�S���Yn��\���`h��������p^��	�O�9X����[mTA���MW���u�'v�jʐ1�_pa3[i< q77�@�`������#L}��(!����b��䦶}�\d��/�i��6t,�m�7�����\���d�jm�f�RƑ����J���(V'�ð3,���!��)W�YR�;�rf>���L��1�:�E{}����3��V��*ؼn�ex�:��M��]}}(� �۔W�����[���2?����  ���Ft�~�h�Rv$^�?;�=�uZm#R:��+�;e��0�[E��e����+T+C���%��B�Ϳ ����]�W�Lz����m|��X�%�)�`�c��-,�U����%bZ�X,��q*TŌ�ng���0kDWyk��X{�b�����%�e�X*$-�[��ry�!;�� : tF^���g�6��6�B��F��e����Y�F��VH�Hˏw�!��1�:w� ��\V��v]-��@pp��`c�N̙�xBr���ܮ^w�=�������8�����uNC�