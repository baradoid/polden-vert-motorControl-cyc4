��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O���WPZ�l�-^ZC�9�juu��`=�t�,{��&�q�^޿��b2	���咎;,���/;{zA��vZq.82s�Y�.׆>�;H>��L�09�JH�q�lV��W��5h�&�|g�-%�_���:�L�6"\�9�v�wo�*��ŭ`�N���E#��#�)Ǹ7��ki�S<#��5@$�tn6'�2���7���o�[���0��,�-U��˥	}Njk�!�����^����S���z�$�TauiEy�iR�E<��2@Jb)��}4�p�#�N6�$n�d��=�M�M8��B��v�R�_���o��X�x�x	�D�%�UJ�J}m��{����4;\!��%'+��&X(�Ҽ�!m� ��=Wϋ3��v��&�:���k���K�o��ل�A�3�ȋ�DNW�ߚSR�E�:����J� ��ҿy1�
NP:��h���2��Cn�HT��M��9��̚�@Z�q�"���	�N���Ɲ�=ĉ���.��!����$��Pntl�-��v`��[���c����L��<!�q���<�[��b��E�O�DX��� ���㾙sj��e1�N\6)a�m��̩I�:#:R��д�z����]L������,�V]�Md<8�pܰ��:���f�r�,8Re3lt�s7t"���lʢ