��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�`���=��5 WkY�:q!���xqr��Vh��d��ikl��L&=�+뼧�=H2~J=*�ʁ܌d�q��q���0>x�qU��q�tҠ��4����x�|���LS`ͮ��zd����C[]�U�����EE71 ���-5����f%�Y��g��k(%;	b��t�UԳS,��n_����|�˜�ck�K�CX�(����]4�!M�_� ;fΌ�K��� g�A�{LD�!��/u�������W������m)�}k��;����W��ѱJR�D�c*#�Y{�2>��Vi�J����H��������Ac��%�:	r��u��q҈��#�_�x��i	Q�C_mka�Id��q��H$��*+*g3QƮ5e8Xk�qr�(�kx���J�0Ƃsc�NF��5��9�9be�2cF��-y?j��u�
l�]����ݷ'��}�{�v�VE�w�& �r�E<{�oТ����Pxq�]�:�wJ���ՠ���эDмU<h�\��.j�Ϡ�<D��y��W*S��
b�v_Lu�9�����;3_���Kʛ}ʾ��_@+�S�T9g�uK¥�oG�1�M$��|��7s�d������1�ܽD|3�&x�NW�s��l@ַ�Lו�R�z1�Nt��}{�ۓ=؉|Q�a�e�dZ%��%�ī;͡��T|�u�_�Ӻ��A�3���
�7މ�h��V������x���/�U�87#ས��T�Sh|�Y�J�Y3J��j������֚���~��BG��[ĽߑH��D�6Ⱥ�Å���ܶ��&fE�X��-�ŋ�V�]z^w��h�#�8��e%B`+�H �7,�� ���@��S(����bi��U����v��
��"y�_���~�?Ä�.�#Q��Ҩ����ܡ��\���in!Өj�b��~�sg�iI�Lm�N�L^��n]�+����!����X�E�~\�Ck�'��r���=�'��Q����Jؙ�M(vҀ>O�"���o�H��5Y���4;��,G%����mGOt��~nd��=�����D�Un�,�2/��)}�ʙ'#� �'�.��;��5�� 7�7�>�+�x!\*��oT8W���]��߸Y�\Y��h��r�,�E l���E�T��q������C�ņOL��!2�-�~b��W�:�u˩!�r��B Q�|(8&3t��(�1!�j ��AY��V��ug#�_���~$����7���S�&��H�Ȇ�V܅������X��dv-��`���i9n�ˑh��>� �r}�.8Z��S��5���&�m�uw��8D��).׍	���r�'&�g���'}�3v�i�L6/;�n�)��)?Ƭ��D<���V���T_=`ۡ����ۇo��DȉO0`m˄�~��/m+W�'0��q�F¢gbzKc��P�}5���2��94|,ǣ�z-^��)V����N����b����?׍7bғ=Й�'�Iv�vl�Y�5R0�)D�?(KaUB�f��-�D�7���9U���8��\k�l0����<GL�������H S������@溘b�>}�o���I�)Z�
T����f;����#�"y�:����DY�O.�L��W�*U�pFe}�q��`������B���9��a}���_�Kʹ|�9� &#�3����j�����V�0�'Rᛡk��W"��,�^�5(�Z�hz����N�bä�5��.$st�wE9�p�붲#��/q)ؾ�R.;F4Nz#qF|YU�|'�9w����N�8w 7)�����@�K�;�B��i��t�}��ik�GÒh膍B���U`9ʒ��vL16�dk��!mEΥl�0��7&4Y�'��5G��?��7������@�Zq~�ʴ�[g�;�ENn���r�gg�j��ڐ�	u����