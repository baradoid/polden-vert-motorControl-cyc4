��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O���kâUP	~NS��d�/�p�I���S.�$�/Z�hOP��� �D����T�#��sR�;qw'�T�}��ʃ�(�(9%�=d��Q�#���� �d����F�A���KN"3$:x�+6�m��C{��VF!��2s���WFQ����Cr���|���!�QN^J^��]��9��&��*���5ݤ��<!.�4���|��sI*���W�ȇ�^H��:��P$HXIe&=��!�~$0vi�&����)�BNZ��;9�h2~]��}���Ŧ��������`����p���Tw���c�p�E��xm$F�j>kh�����$	��к\��|��i(�Wky>�2B׍�W+�Ŏ�G���~�-�a�l��*�6[`}	���io�[EϦ5����s�EN�hC��Dǒ����b4��T�