��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��[��&�f�u읪|�9}*����Y:T����Y����,1 0��F�1�0պ�,�9J���(�S)���M_�0�n��[Lܲ�}T�t�/jv���*�9�6����@�.����R������ŝ�]�?�K�%É��&�6���k��.Po�S[���֯�=S�&	���*f4�����<��&'Nj��a�
%��x�Eo���;<D�H��\�#|�� �9PK�]����T��y'.q
D�Kk����E�Co5������~w�[L�C���F�U�O�!���������>q.�;���}�}t�vmz>"��dn���R���7������ѡ��+������%�|�sp���ah����m��h��j޸=t
�3j��_'@L$W��+�NK����&2����ơL۪�
�7�(��7n�w��`�x�W �-�gx����p���N�f	�7�~��|C]�}�X��ϰ�.b�*�l.;���-	��Z�ĥ�Tɱ�٢�L���I� �r��b��k�&�zi�k��I��5�ӧ��W&>1����qR
�<�m߸��Jf{�8���m�F�"PY�����Φ�����Aٖ�r��ܝ�}`��I��ԡC1�,��~��m�}�IӍ��7K��餆�a�Q�檽�k�P��W�E�6��1D*�Q��O��}��ؒ&S���8-KЬ6u� q��ᒫ��ʺ��GLf`%��������R�4Ϣ���7Րk~���#�*�����Ӈ��:E��L��}�I�L�����͞��}PA��N;��"$GdF�/��.�gm�$Z. +�}2�t-�s2�XÂ��4��/Tet(�{z�)Kr+��#�*� 㷌MoV{����Az��jW�5wl�9��4��#��,���u�����cc��9G�VlE��j^�U��J%��24�Ol>����1�9q�!Y��� �s��L�LdH�X�F���	3�u!�FJX���{�e�b���Kc/��nx_8�G�qt]F	�%�h�ۿ"�[��7����}�A͖�/����3���藍�%�e83�Ƨ�Q�e��r	����R9�������@/GX�F���I ���E���@#Je��LB�(VB>΢ �2�����`�8}D8�U�13�=���~�X�"4ú,XrT]�����7[�g��쪑.Ն
����ϣ�V�<�;Se�[d�|�IfK؂J��;�o��AǷ��D٦�.˝�/	��Ƙ��JW$o�e.��o�Ȓ����?��m�)k>Ȥn�gy���K��5
��d���N�����Sh�A���Kە��
tK5	N;m�h����|`���ƞ�.��4gm�/Py�����w��������f��	�SM2��-���6@	���/a���N�� 7N#s��z���wC ��[a��{ ��3YJ���~t�y��'	��{At���U�YJT`����z��_���ME���+�ە�� k���~�Ѳ��?~�ľ����(�xl~(L*�L��NY�4�{�qr����c:�,�8�4����Nb�2*ψ���٥.jÑV�Y�Eu����-�
6I�j�J^& �s�S������M�0`��b�ô����K�Rn�2VQ�q�@i���GП�p��]Y����:��[_���r����w�e��;�<5p��#h�����_��*_S'g-�ߨ�?��͞vW�׫O��:U�5�f�K�t����=�m�?�cJ�c��XpD����FO�0RR_`��sf��^Qw�RĖ����0��oqCM��nb0����eѿ9�6_=�Gw��H ���9N�+�6���XM��ǀ!�~qG�ZЅi��x��5����8�ת�p��"O5�0_�>ܗLbT�(�.a�Ep�����&m��%<]?��m����Ƭ~w![����:2�G�~��ϗbK�~"��i'�oW�z���7�+����p�f�։ɥVd��֬�O�j��.���a�5D��b���	>�̃Pv�W��B�X=�2e{��8�g�#P��7\�����yZ8�)sk60�u������A��Ji-���_g�o�2.�8o��MlY�eU�q����K�#��j�jkP���c�ks[���uG���n��S�L�iy��kG��R7����ٺ,���&5��c5��W����+�����
�j��m��.*��S�cn�I�g�yH5	O�3��QY�*�"8~�+J��D�(���Z�ꑆj�(Y0���f�{I@j��u��R��j~p�!L��ǟ��l�r<�ynJ�E ڙ��X>wx���EV@i�+fd�y1%2�[�8)�7�2q:'��D�2Σ�}%�h�
�[�O�ؼ*�-�o�d�OQ���Ż�b_n�9�� _(��u͏�����Koʗ2$������z ���0(@�w��7���+���G�,s�0����� ͠�K˾Y0����NY�I�*�w�.�F�_�Q�֔;�2	9RV�@�!�F��YTP$3��S����;/�	Z�e���\`��yo�z|�W(6�v����T�$ �Th�~G��
ї
3��|�T��k����ʞI���7�/����̌��g�eP)>Bp����[��ӫ���ˀ�]��F�3ۃ_r�JmJE�%h���$��M�:W\H�g�.�Mm��Y�ӑ$�p���9/�o�f�짆��Y�#��M���Y�E��y��!rx����X���:�㘈��/b��ROj��� #M�0{�|��@��4��4��\n�Χ ��aʄ��~���^4TRt/��<U�;=�6��襋b���{���j���[�V]�k����%�
¨��F���/��� �1@��8�ݍ�%i���A��˱����qsj��,@s����ǲ��^y���s��}��{B��H�Eö�vK;.,�̓ԙd*�no���b�eݏc����P#�ũ�#�+���H�UCp�dN�Om��6�8/���BJ���������d�Yu��(3��Ui�W�e��HH�)x�FJ������9�W���[��>q��*_B�M�Q$���C�&uy�)DG�=��\\��^N�
^��w�!���A���@~;��]��~�9֍�n��g��c�O��m�+?���CC+�l�'��U>O��rl�vH����#��/=��F���������2F�E'	�@'�r�]_��@��o�&.��b�p�7��
��֞��=�L%�Mͭ=��xڣJ��#��/5e���qE��w#��37�A���z�SS���"�\5u�?�y�[/6o;.қ�۴��K10���,#dV�l�n�kX�tҧ�I(g��b���1�4���7<�a�.����"N� 	k���=�a��_����E��|�?������&je��j��%r]������8ePYb���~��P됲�����{�
禨��h�!�PWt�\�9�A�ݨ�"����Vm�E{����@�c�Id��x��bu��ڎ�K cP\�[h���%_��� ��1�;��A��>+ni�mӍT���B�?S���D�o>�:ڮ����[����x�s���Y����}��wSF�2-������(�1gb?�3�o�P��EH�|��ۧ������A�H�8""����!�w��N��9����l���q�1�q�OX_v"�v�"��1�oZ|�檦��a��A�BCq�X��_ل��+!�} �o	����l��כ����6J�m�?��4]ѭb߽�.�8�
b9�Iop�&�)�;���d��A%�"ʽ"�/�ㄉr���T��	�s��f}!�L|~�L�\��U����W����`���\��To3���~v,[<| Ĺ����+	��q����S6����(iT�/Ls�a12ĕ��|�/�+���4�?D����~.�C�,�c����=��j�I@�n)�}ԋr��u|���l�HJ�콂V�m4�D��؀��~� �'��$��Q~��������M�ׯS%̿)��-���|��roCu�1�Sv�����a����!T�h52��n,�a�AY��֫��|��+HP+�9�^��ǒNSـ%��e��UW3e
�JS����+�R��y�|��J���%h��֌V������������w(n�,�d���f��ځ���K�4?��XA��Nҽ���N�g�
WE��v��#�x f�|D����{�Fʏ	B��_� �kEؚ!�^�T�}D�?*���)��X�jNT�2��|� �;&4"Cy�r��uT�xxwPq�����Ȣ�܋���X"�Æ�A
��"@=P�����2n=/������r��E�&���x`��F3N���b���
Nż;h�u�ݏy�.��B���?���y#��>�س�M0�w4�F��--���e�.>Y�'!i[�>N��]Թ�Z��s�>��5bŦ̬�,g�`�{q��9#��g{Ԃ�����ɗ^���3�_�Ɓ~�xߝ�����_h<�:�1��)���g�$5�'d���u"K��$/k?�_{b���f�T>��7P�S�+�e����2�p��3�i
*8Ƥ���͡�|7�q����U���N?�������n�ޯ����F\Ń����AzF5z�)k����~&t��u�շs�����x[dD�2;3�B�0,mEkG�:>{�m���u�����&�QW��!'��<��РK96�+e$O;DAM=����\��B��sf�@�=Y}K��t��8���e�-��E�H2����-�=�;k���W��6�/��al
�÷�O��."�Y���K|�ay�~��.q1[Ű�$�@��r��<T��fb�K���U���D�C�$�I)�D����� |��p�O���������9 /`Bj�täp��3r"(c�y��&���:�2���.���R���k�挧��WKƤ��uM B�_�g�����w��.�i9�%�}�U@$o���~3 e��>;� �h�(����V��������b%I�4Uh�	��wG��@}��9�����Uw�|0�YFfse���<!�>�Y�h��P�����/�������`�J
��j��fr��$�EV�*�{��4�~�q,3iߔÇ�\5�n�����r�<4�����������ɍ)����Z����՚��b ���ڥ�c$fR�٩K;lD���w@;�H�2'b^��:�D�యt1^�Vo|Gv7o��!��俐��}�}G��_��(�2�;�M|��,��"���e-|�ŅN�3.*�����J��,�|�;�`ٲ�9�9�D�6���|=A!g��l�Q��R.���W*�����K�H�Hm�=j�����_K�G�����"�n�{yv�������^��(Y6ć�s��3����rU#�dCJV��G8/���s� �.L��]�F��bN��iFI
&���O,8�A9KvMBFpt���MN�5�f �CX��o�F+YdҚm��e��]��k�^F�w����q�@dX|�"�����C�܍˞i�ϊ �H��5D��G�fڬK�;�fJ�˧x��E���R�%��+D�爞i�����v&%ה�"ֆK(��DW��=�s�&��|�$�*o)�7�O#���ȃ��\MI�'j�I�1���rPƲ�a�a
����Km�/�s�6�)7�\���R5��+�Y�TL$�.u�>�A�tB��o��y�FGr��;<I�Fq��vK��*�"j��ֶ}7�yƒ�#��+E�T��	�te}�_�u#6�u� �L�_m���%�N���4A���B;ç��� ��D�~�C�����*���vϓ��V��й|4��Cg? U~�C�S�~`�T�AN�!v]�&	O f��"G����lJ�t~��*�|쐔�8!%�7�/��j�>2�k���N�8�C�SZѾBi^�s�(�l�c���gIh0�������dh�D��2fV�ʖ��0;�����>��jQ�[d�ܤ��q�bތ7�$��m�u�ӣ�9�Pl����W�A+ɞ������h�Xd�l�C��΁m��J�}��j�����Y���-� c�e񧪓��>ߝ���U�V@_��m�q�(�4� h��u�|��ؑ��C�`O����EA�-?��JM	x�R'����^σ[I��g��U镩e�=ۯ��xN���KO��;y�]�9��7�`k}��ay��q�뒡��@!y٠�/��8��Ez埓�/�Jk�������`�+��vӞjN�(n�O�;ҙ��&	�*�>:�P�Imo�cg��Z<�a���Ʀ=F�!��% �[�����EM�O9�}�~�^�K��I=���?\Xd�$��
9�S�F��b�MH��<B��mx R���˧+���[��������Xb?�8���m+�L���$#��P4������tJ [≳�w����#p�u���QZ�y�VW��w��Ҽ/
r������8�M�"ܾ��B8�R~�kV�]�j���d�@��WB0�L<���=i���I׹�TUM糕�I�A����k�@�@�D"wd�i�|�
�ǳAC��
3h�$���k�*5�sˡ*�ӦK��O�o!��N^��ɛ�{�h78/)�tʛ���5Վ\��hz�B5��=�W�s�]~�q��#?*`�"<�� ��?���X���ÅQ����#�qLд�]���7��s����|���?��
i��w�j5��i�+�����oވ�yE0��#W,�x�~�E-/��F�~�UpJ����k�|��RϬw��R���6~�)��,Loo�8�у*�:�/)�B�{#:���]��D��֑Y�"���u436Ԋ�=�5mRB���\	��U�F�/�|���w���cr4��6���qޢ�i
���9������������*h"9/�5�^���\h��a��;��}�"�.����)����TU���t0��;-�z���ߞ= k\J6����T{���<��	YK�GubPU��Gd}O(/���!�zSA��O-���Y���,q�&sv󗗻�hT�SR8�p����ꍒ?<&p�jUm�.�i�Y�O)����3J$&�h(� mt�N����_)����O%�Ha�XTO�K��m�˖���<Uw�ܹ���e(C�W>�;�S�]�9nB����g��:k�l�j�̵J�%%V�$5Nz�v��S v�U��K���m��St� ������q�ùÌ�ՙ�@�;�w�	L��^��䞼6y(����-�*���x�����������*���d%*�P�P��z�q��ĳ)�������2�CG��ʣ���rl�,x�l�8�7�� g֨�׃+�d3�v$T�� A-h��,�pd�џ�C�\ʊ��}zKk��=��f
�9�Ɔ[F��ZJ��ѪC�����!���K�頞�jb4�ک�l����S =h����h&�s��U��Ƽ�l���߼oT���+��|��)�t�S���V��U��6\�d�UG�>�sE�Ի�����J��<͙ �1╾��
i��`I.��	�����U��2j�sjUx���j{��1j�6��;,6$�A੊&\^�3�����Ú���9�y��g�͆O(�����NN�z�S��>p���������T�{�?�����ț�?-�̒>�~��f���Ƣ�:�t�Z�;�t����[���a&�F-n ����
%�/���C����!�;����և]�e�
�P#��B�p����U�M��G��,$[��Vb�<崑e�@�Vwuԙ����{�_��<`�jJ��P.��j�C+�aA�~s����|}z^Z��l�=lׄ��
G�E��q�Ä��l�͡/�d�wYb��Z�D����X@r��[�2fu�Ѭo~���ġ`�K�r��W�á���ӆ,=#,�F~w]�0�^=(��5�j�G�oq�����t��8���_4�������a��	ؒbb/��x"p���n�-L�G`Ң�i��K'\B�R�hs$[��X{T��0��t��J�nE1"Sdn�����\$��[���<B������z:D��]DH9���2�z���7�M����u�{R���3&�p�PB��8�a�����&��.q�)lr���?�[PwkƃV' ����� ��%�/�O�d����(�xf`�щ�V�â�L?��c/�j��Yq�OZ�
�PtoG������3��H�6Sy�%�����|�\�wĵ��%�u� ��cy.=�E��T3�0��^:�����Ǳz���꘼-Ȏ���<��]�X��t����,���)~Ti��p���-��{�>��LZ�	7D��C�;p�.�"Z��cM�(�Gv��X����{f:����R/\p]�;g�Ss���b�4z͢�J���ă�1K:*Q㼰�F=��K̂�1ַ;�T+��GB��nS&��j۞'���_��Yr�O!��9$���
���8B��ld��6�.E���ryܤ&���� ��� "s��WM�� ���^������`&�u�eK2�����C����ma����&��/���ǂ̎r�k����2�,�ő�O�sw�D��G-ozjj~'���d0���q��&�ʔbS��D��M�-�^�PN�"9���pa��]9��*�V���6M桝�n��+�����N�ߧQL�:�h��g���XM�6���
8�bZt%�߹�#�R��$���D�w��p���;�����C��2����f�;brd�k����k�	׫m���Nk!f���U%�q*��ҷQ����;ϣ�A�r�lU�fT����Y�)Rz�Z]rj
K'���Ʋګ�.��XlރWђg�5��=�܌�]�'���J��a�kʻD�fE*~�h���u��\���7��^���e�]�P�J��TV)�U-qu�z2��sK;2bp�-�D�K$Z���9��X��Z��S����8��?gz�`�OǛwˏ�{N��\�����;���KUP�%��0�U�T�M�zb�jh�r�-oO�2
`M�k�&����ɛm�"Jr�<|W!n\T�����o��~mi%�_�^�m�k^�0�9B��P�}�d��&/mv���R+�IW�4n�`B��ʽg{�3H�Gk���H	!���U�E&K��o�[���7�"sO�츦"ǖ����!���Pt�hD�~�E?($��q �pY�;_`n�g�: �&����M�3�/!cʯvB�9ޔ� U�5q�~�����\�'XOp��9lSw���A0��L<b����C�~6�;
8�5��o�b�x����1�7��U�<�;(��|~FM}�aF���p��)���hE�g��9��N�3�Rd��~�<�~�B��!�{���?�lE��
�|Ԭ�	�(��ʂ����Ů�A��0F��x��0фW�`^,��;�����?N�:k$��<Ŀ�����4N�`�Zr%�g��!z٘��tTb�ps16y+P�߀㄄N�����x��I�A���h�����	r�Zf� ��?z�2�8J��������� ϼ�n�&�l�{0�
L�3�si`�-X]M�+%�co>Al.t���L�]�7�:�2XI|�	��ެgdIH��l�Y���6��\�<\���!��&0�,�� �>�9&��E��z͑Hq����Eާ�F��\�pd����]�t߉O�C��� �*�ͱ_1��-�u�����m�}^I���w��I�^Tm��t6Lq0|"f���Zg�N]�3b��g{�Sy�P�cwN%�1Y�U)IxA���W����t��+����#���A�q�Y�W�������wg�k�f�ʜ����Z�]��*H�r26��,�&�}���5d,@·�L#��n2k�$H��;���J�����9^fq��_l W	<�%m�0`�8�a�3��]���_P�7_�;@�9�@��E�N�>� �`��0p�T�/)��:���`g�&n{l��a-�O͊C�vvT����r�N�A:|��2�}�9�b��B����T�F�0�	!(���@N�1l()i�$�Yczts�.OeF3�v��Dиl��ɤ�d�-�!=��+�E�l~��T'�m�S���
��,9D�1`��q@K޵u�k'z8�F�jɠޝE$q7ܩ���t��5��!�E����xف���	�O�ƦVժt$@���N)���	�J>,�5�Og�\Z��_�j�$0?6��Kj�2�D�i`��������)rJ�����k���55~����r��,�]�u�ZB���J�'�Վ(w�=�d��2a6�@��� $9S���\�د��X4,c�]ur��}YX1b<i�sD�PDW�%������z��ϻ_~�S5��=����k϶�V���)�k� ^��%�� ��N��8�ñ���0|�q݊�3��|���&.�C��K��7���#�yj�Z�w��V��}^L��E� 9��܌ ����Y��y�ĳ�D��F���X�4���َ�'<�mWz��37{�ߪ�3��	���xyM�jV��׿Bc�Ӵ!�8� ����8�g6���:��>��o<���yc��NbDBl����=�u����7UaU*�,xL�p��O�NW��d�c%z�=�$��q9=Vu�X��w�ר���
g!�j���{ȥ��1�v������X�r��;>.G��C7��F0��-k	nf)'ufDU��f�敐:μ�؂
S���#L���4r����A��f�`�hTw���H�*eb�h%��u���:��I�Ǥ�z����iQB��~RHZ� қ���y����4����V|
iy�����ȑ�>I�[�%V�P����N��Z����Zw�Ȥ"#�)h�r$.�%@��$�v�3j[�(��Dl��u[n�N�X�2cQ�&|�m��
l�aUm�`�\͞�6"�#�/\���H��C�a����Su�^�l18k~�z˄�y{�r�0�ѝ �{$���aV&��m�B��8�O�w�?۴�j�T8���o�ȣc���#$S��z�HE�-��������eWV��:hW]����hZ���~m�l��L;e�Z��M��f�#�Y�7_����`W:��1��6a��nÜnH��*��X>�ܔ������õآ?,���B��g�����U��(�9۹�6�'l�ae* Ƣ���{�J0^��C��H�����w�x	=�t@���xn�9�֓�+��[��@b����"N�"�dWg׶�Y|�v�]�Iӄ�Kt1�!�"�W������8 ��I~^Ǹ$�d0'�,[�6��S���' xx3!�ѻ�ڢA���|�Yݨ����t�tPy��ؓҭQ�O�R`` ��٢��\,� �V'��q�
[S�E�q�!X�5Оp���V�7��T�S��~m�"�z�-7��ņp0ƏM%w ���Քa�[�]�W��6�L�V��w��/��p�b�}�f,8pF�8��nh�����:t��������������$�[�H�\X������*�l	�I���M�D���A޶j^K������q�+o"'	z���P�U�ZЯ��b:��%�I