��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�=l��!ӻIA&{7��m�cpԼQ�J���Yk��6x���6	���T*�*x��ǿ�Y��p�l�s��RG�\��@��o�G��d�ZM����b���Ѝ�ԃ�V!O��ÿ���Q�����ʖ�	�B�G�|m:��[�� K_s��<kZ��>�'5����C�}�cj��ϭ���*�V����t��7�����05��b�GH�c�f���&�iS!IӲdE�k��B��z����n$���T���T�#�o�L�y���5Q�c�bTt�%�����]��c�!�Pu���"���_�*�R`�V������e�:�w�RML�@o�B�#s�'���7	ϥYta����'���n X1�L{y
�K�IT^�A���5�J٩�1���&E�,S�(]�6^ Ib�j�� �kr��K��r�M-e�����C4�����/8~���s<Do���+y���U�~	"Z�mK:�{�/ ���"�R��=�}�x�!k/z;��%A%�HH���T�[ ]~LAf]JN��v���"IU�J-��n�)�{���� ��H���-L�>;?�����6)jc<w��1�*�o P��Pt�MI�˦��:�:7��7�̋���.H�DU��TKH<e*��:ޛV\�v(�HF�̓��P����(���2$6`�tg���H\�T!��R?�JY�<6�fY:)��c�A�:����_ڡ��R
� ��N0�v��h�����Q]s�����y�Ӓ�I�E�J�*Q����\��:ow˹u���͸;3��: ��1
����P�M���|#&�s��{����jp	�^�.��r�E�+(b�bs��z�KD-WX�^˂�04�qxT@��Dm���i�)T��'�H�3��!�-��{�̨�mL�6�_L��Au�L �v3l�|]y(�	�#eX�5%O	:I��>*��&��|뱂�leT�}�͉��2p'_��.y8֖���'�n#ꨜppy�%hu\��qdѝ�4��)�˨{�(q��6r�܋SM�&|�m���d��`Ou��`��u�.������~���|���=}K�E�ӄ�����@��n'pcD�v��&��S�=����f��#Ɂ��U��?n�BJ`O�ơj������Ab=�Zm�u!|M����ҍl���Σ�� �wP��]�*��/B���6�~K��9. �/�t_I��p�r�ՅC�4.�@��:�O�x�t9χ�u���>��2��&X,����#�̱47�qe�j�K�ܭ�#*�n~M��]��F�ZrIݧ"�t�j 1'���w���G��/��sDQ�2��^/*S~�����f8���J���8����4ć!
�hc_��e7�3�'IҙV�Q�{�$+0���|�=�$���.�ͱ����Ђ��T
I�̉�[l_+��Q�L��4��[7��Џ���Qeuf��	����	wg�^{� ����_���>D|��[�%��w ��
8��ٜ��r��X����r.��e��N�_2����Z�I�2�m���g���������o�*�ԏ�r�0Y�R�P�g��x���+:[5��J�� ���B~�2_;:�o=�����P�C��Z~��Ϧ`a��M�
O�#�����S�0��(�Z��WEA��<I&��R�fT'}#B4�&J���!qg�v�O7^qR��݇@�?��'�y�4%��Ü���%-*�L��L�f-���O�F����3h�y��E̟-�Z5{�����~��bBʉ���� �"�ht���\;'Xr&ݜ�D����1~SN��C���gJ�T�L�_+R3����\`��~�y�{�'@������(�*n.�),�H��2�X(n�6sC0�.���wh�1xa��zx�50� *1�|,^��N���<���%_h��Y�X	�7�xbq�ӪA����$+=���߫�?����/z�y~���77�����or���@��Au��L���@d����G�{�iϒ�8Ż2R)�N����9�St���$M�ܧ�X�:Zٓ���&���&�,[C��l���I�ܭ�6��h:�c�y��H���nW�tʲ`����(�+��b&N�~� ��\D}�|&	'�#PZ�)4ʑ���J����)4���<S�j�l�b�D������O#��3����a����MC�&�2,x��h���,� =HDM��,���90�2��� ��c��I��7A}U��}��&�n�U.�����D��g��LuD�9"�.�J������$̐�b���y�m�ɶ�:�L��� 򱿄�*~���>�t�~(J�C�2J�����SHD,:R��NBT�#w�僼�i�{�NY�<�K��-X�{w.J7��T�<�C��k�N�����F�Ĩ�AWe�T��-�F�˶{���4J,�`5<\O�+�ZL���^���oE�H���4I�r�`YJ����P���o%fF-a�{�/�=�G��iL;w��+�#�� S�:��\��ڪ�Qו�!�?��;����_��v
ʉ��(	�l�-��R��QdV�%�9"}.��ݠ	BP�Q?��z䣽�ʠ�< �b�����;�$�!#���UN�����1���k��ٽ$Դk9n���`�,Ws�Gꔢ��J�;�(�D���q��B�ÇQ0!/J�/:	b��7ҁ���"@�@�;��o

?�lͥ�̓���0�,b���%��߅�U<)V:��G]����T�1a�A�|ȱ1��Б7��h3IuQ��a�
{뀁�%�ó*���4HQ	�����'�2s�2׷�����aW!c�Ȉ��.
K�g��
��@��
�~�篽���>G,@Rd��3:x_��3q�nI���H�F�P�p�~�s��7���%Ƨ-u���Bw;pcv��殌C�����v�EK!��C3�%�f0(1���;g�)���S�K����g<��(����FU�G��z�������UQF�������\��b��x�M��H�*!+�diǖ��0���7o��gU�����,��x��(�V[>d�1���q�����]Y�e����t��&��4�BV�^����� J�E����[���pp�l�g���)�J,�6�^�"W����\{�M�7�`���e�^���|"DG,9���eI\������~HV
�᥃Ce�RT�g�м�Ү�2f�㻊�_�T��~���^�Ρ9�
�-���sЮϮ�
�7x����"I�9��;nY�R�B�}+�*�XbԽ����-Q�o��i�4ӛ3۲u��.��q�J��2-~I<i-�ߜI�DI'5>h2Z/Vv5~6Xͬ���k�EA��Ȣ _��
�)�w~�a�n#.$�й)�1ίlX��c�n~������@����c�W~U$1��X��
�b�GD#�g"�����#��Ja�9�����j�8	��#AfO��I�u�Y�k�Ml`A����9�t�ώ���#N^��w��F�M���8���#�8+~���-� 19<�b���Zږ;6V��%��A��8�sK�AaY&ے�& uSc�q�W՝�<6��i��*ßр:������6�o{��s�Ѷ�����ah���beq?�1�Cd����9gjޛR���+����UU)V✏R�-9J��E9ouu:'w�\0��y�Q���}��y�P�@$��ƭ9�	�~>���e�gJ� 	�ۭk���p�k�_(~]���C�/<䉐TkKALs���E܅O��+�qF��"�z4�����W�����:�pe۝bQ/�N����!�D{�vnj#�7x�3�T?'o�{�d;���+>>�[7^�[S��0o��V�_]k�&\�1^�8;�\G����̪K�q��o0N��Z��?�5)��<t�PyA�t���񳵡��h�:�&=�6XS�	���'��=�Y\����^Y�����(1��ҏ���ɫ�옿�����'nv�r~j{�=9�Ps���-u�(�YD@�E��*�
t�O���O%���s����`�jU�(#�g\�)1���� Ֆ���v�)�L�-*:&Ph��Ո}F�I�P��bH�r�*��6��(��ۘ��l
�i9S	���,S��v?��(��������}��^��U駃�Y�Ӂ<9d�c(��xd�j�2�IJ��b_��ģ�oh�
�5dm�P�Q����6����v���kH��#���2�q��z��.��hq����GB�	���R_�g
Ǜ��rS�cw٬��jۢ�e Ot% VqT]�(���������*��-�d��bs�(G�g��T��">s��kyT�H�v�8$�ƽ]�s#�;��ڡ#<�{��f���Y9TK���������	ݪ�
o��Y��? �|�!��
,mR�����1!y���6\�(�඀Lo�ĥ�apЈ����ӂI|��;EI��˘n�����:4N[v|	�G�?v�� �����}� 3���fpظ�"���;�tM4�\.ϧWE�W��2�w�p��p�֞x;6�D�t'����JAw�ǬQ��-��\��5޺6����h:�!��wD�-�b�]	��ˋ����������?�xN�`��Z��t��@��0FƮ�b ����D�b��+QE &3��\,x@H� ���A~2��I	�b�d]
l���b�>լA�=�FRt�@J�z �,��)� cJsK^3�F�� �Щ���-e��ͅY+W0?���Q_㇖��* W3���I�g��<µ�<9�"u��?���t�S;GPI�Χ�m��pWYm�^�%�(�݀t7��{;i�ݙffm4?N�sI�y��P���r��+m���귕|L
b�q��=��k���_��/m�Ф��7[z��w��N�er�2��6�Z؀�9���4�+N@O�4w��<8�Y~��Wh���_�V4?@F��&p���t�o$|��Fs�#�2�A���W:�6�)��ѴRO��lO������8� R��%5����1-�\B$��(q{���4�"��Ҕ��(y'�2��`�����m��F^J�(闎1�|��jk�L���*�.-���J���ۀZ�E6d� �u�'� ��1��9 d���l�x�BÒG���ѧ� ����M%e�sB�Ă���;�bRN���Cflk��H��q_��ϸ!=����BfY^{��9k#�B�G��|,�`)��1���;+p�Xnj�>"�+��T�9#�� ]�Z^*:��$��$�y��-�f�)Z{Г�����s�6�ҲuXh΀n���=��9o�����xk"8pQ� � ��g��4��f��� LƻO�T���� ����n����n2NB�ֺ��a�2ZV���=�ȖQ����Y���` ��S�7J��,`4�T�GT�$q��3��������@�mҜ*J8���`�Ԩ�:�Tn�H�ܗy��dZa��<?^�+�ѳD��6**a��$��C��?�%3:���������dqx,C7���m�8�$Ə��ߩF���ͤ�M/G7#����C�M5TF����B
�sn)�W����X��jqY�i���yX{���c�A�KD��I@`��a�ߧ�a9N�G���\��L��=l�7�?g5�8�s0O.��`�|>�'K:����m|��YgD7������PhK�������Sx�~�x��E_���)ݶIoy�]����C��t��-e��KA�uP���������IVh.���A�Vs�6�������u��w&�:7���mIn]��}��;ǀ#�$[4y�d6���7�$�35-�m��;V��|2�� ���u��Vg��ְ,-;�X�Z}Ԉn'�3�D�8�ʁT�3 ��i�|չ�k�q���&V�|!$�ξ>�ɗ���^�X�g� �9�[�Q��dZ��B$����^#��h�,cw}h��'��23�i����xM�b���]�����,�-ذ�Z���e���S�Q(uy"B�U)���8>��+#�����T>���k��7/3�Ԧ_��k��n���"�\�Zy�eZv���Ic4��x`�"�z؅a��@��.w��]�����֯)�������@'�����!��"�Z����wn\j���'p�I���Ґ�L�jIJ�Nv��Yzщ�[��%� {�j=�fr��ʕ=i��K�EM�!T.wl��'�F��k�2���<�E�1�oL���n1�b���;mP��[�X.4�D��(?Cǒ:�k~<�ٵ���??�V6��yB2zّ���ޜ��	a���O�����M�hI�����\.��`Mv���A�A�G��6�@Yqn���m����Uӯ���]+�d�zp�ݜ!cU���j5�p�D��6@�t�s��z��yZ;1j�J�.�����L�T�Ȏe��C�1�H�9��k}i��A+N�Ȧ�ql�^�F�R��q��J������,�N����x�E���C�
P�6��'�K
'v>��6�/�S�a�q{A�ɒdXXfi�ܕ�<�����:bn�1-�G����ܮrc��ʖQ��Q�^g���x���-<mBp����o�����-��m���M'���Ʃ����&�vE����`�ƾt�	M�#�-�$��ַ "G�wEna��M()h_A���u�N��v�6r��z���k�I	�*��vZa�iX���� �S���<�Mr 	�{⨻�ǎ�	���l��UgHZ�e�h%_N�>^i�;�[�V��՟��`���6�#�c��Ľ�W?)١�v�|9��q�x<F�Z��ٚ�����lWnih3Tּ*t2����M�������,��&0>�O�A�TS��	�騤,6�Z���Y?V���[�E`����� P-�ZM�_�泊�=�k�@�&�WN3p�[��q����N�F�˰>W��O�vu�,��<e���dκ��=ʜbH�$���F=�g6Y�8��O��ZX-��U�EX�(:�G��e�?/��lÿw,�:�2�ѣ#����5�w
!ڪζ��6 �S#I#p�w�o���G���[_����7y9�(�c��SW?���~���h�L�|ܗ�@o�PV��#d��>��������eG}rg'�_Xi��4wS;]-mD5H�����/xp�����5�B��l�Z8<�8�i� B����u�W�X�j�fA��jO�D�&�ӻ�rK@�[���$qqd�����矸~
aX�Z�2ī|+�,:��ã�p]��O�N.Xa����付��9�bDV��jE-����{��^dhp��\8�I{F:���#p�a[@y���z�9�p�a�,V��&�r,mn "��Z�fQ�!`�$�
Z�ԅ.Z�A�є�LHd��j����� ,Z�e�5�ʋ��x�,�����&7�}gJ��?���0��)m2v����r�/_���y��K�0{��md�z)z��2#�{v������>(��'5�}�t�v«)b\��}�Q�r+�rj���ݵ�J[�[\���H��6Їb�X��dB��6'F�ʆ��W��5�1x��`q��������L����}0c��$����V,R�a�b��8�³�絏�r����i+]�wn/��[��)x�Z�90I�/0�񲲃�����^V=��G�"�@Kw�13���.��mcU���e_֜+Ne�*>h#ۂH0�V��!��%7�e?)�s���d�b-������� ���2^]v�~��7ƹ�%W��}i��17Ik�����U�� �ŉ��@C*�B�-�F��H�2_ZA&$�.�jB�I�>+М)�&gp�\�=����Z���)�d-"�H>���Ø�w�c
�'|�� ��#<4��mOv63p���S܅��P:%�~�_uO��@2���+$s��v@�����e5̽Xf��b�s���^$a���2n>�������a$yktMQ�!�)��T3;�71�a����!��D+���dX�_S