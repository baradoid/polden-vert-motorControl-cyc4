��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�=l��!ӻIA&{7�Q����'v"_61�'��l�1��P�����s�b��x(�yϔ�v�I��ǣ��?�����w�n���!h���,�e�X\`�����}'�9�}��n�J�n������X�z��s�'3p��4�y�;�7ӧ���M���֯\}�%pIƄPU�Nӄ]���߭�J�%����Kl�?��=�M:�BX]Á���B�9͆���|CA����n�&�^w���2=�Fzb�__�In|1�<�~`5�ˇ<gFu��r���q9�i�rEG���N|��\�z@�W���B�S-w׈}�O���.�@��|��9ȋ�.O�[����7to��>Z'Q/��V�_��zy؄�X,�.�	\t��� ���^v)���]����=��U�+�%P�/�3΀����Y9�Vͳ%Ȯ	z�,z|��!%�P����kv��h���i�r)u�m��?�
�	xH��� ��N��ṓL��"��3���Z�'T1I�mC���0�:�c�����ˤv�P����R����&�xd&���Xb)����Bc���.!�5&(Hr�,���kE�W�䛚��Y;�^�J��V�V�%h��?CH�G��w�m򥐴+`�߫�'?�`�s:���(�%�@	ɵ/���>����z�L�ύ����	���x�ݡK�`�(�^��ӎ�Dx%��{<TLo�Y�K	�~���"nWT��AL��b6
�W�~߁�b88�W�`�RM񻿾P���!��������b�)��DU{�\�|(�\�Z�:K��=�"�F�=�02��)�w�����&3o��Ue��,|Q�\A���<�7��Z���[nL����隺'�X�w��g�+�� "�6�� ߨs�9е�u`��ߕ^��e�A���6�JT
�^�5" � ���z�m���}�b2�1ռ����<���0�����懚�0Y�P����5C����f/03������f�Z�%�m=��sbP�<�%��Ji�>�R�>ǹ�s�"&�&�,]�4đO��k��3��,�ւ�����[���'��-Z���m1�d�'���|�J��j�ѧJYS�ԛ����4�$r��M�֓��Fɥ��^RW�/��4k{��XK�I�x]����"������6�ߓ�	�es4*���b?�頢wd�1�ٔ����h��rED?����.�1�KH}�8U�{��������$ms� k���%E䅚�9"j��3f�D�̡tqN��L�:`S�6�rz�P�l�R	�(��pQ��ˢDTѕ:�Y:����*NCs_�nd��^����Lk�eԦ��~LɃc��\����y�[�39��^�֐q���&94�z֏Y��N�:$�to���^"HՒxC�G�YQ�����o�&X�*����J>���x�������g�i8hp�x�Y���W{u[&���R�m�A��\�W����:V��qP�Q俹;[�^�Y��y���:@#S7�!oN �pl�)��ꑝn��
�b�ǯ-�	k���v�!V 6��rv�����[N/c�Cӓ�������,�L̑x��{�QtC��	ٲ�~B�{>	���%�U���\	(Q^�����ʹ_��"�{�����WĨ�s���<E�)��*���B��(��Gs8zD��t]�����2�  ����y���;��� �*����K=e��憸x!�|�v�v?:Ӭ�fD��L�_\��xu�C�cr�6��:B@���1��%<7�n�!YqTVʤތm[>\6��P�s�;��7��������s7F��	)�������?��`��P+n̛G�-�I�U�����~0����W�*��ޢ�m�6N���J}Ѝ��P:�t�OA���7�rMM���:zے���P�E�蓊DM	��VT�@F�5�����)�t@W�����L�MX�XA��p`ē�>�~H�t���،&FJ�dO��=B�ua�r3�c|�^<��a6���^ ���!v]�SÎ޲��N*T@4��!�1U�Yqi�K*K�2��L��]	C\�g��F�� ��3��j���T�J5��"w�@�M����K>��j��V�씷#UQM{JSz䥮�Z��]�3��[��|^���#�mT�"RX��O8^U/��
���`FL�J*Ο4'D�S�����ӳ~$�|�USݥ<ܖ>����T1
�P���B�x=����f�y���|W�u�s�������F\x�vC2M=@\s�]�IΙ>�Z���&K`�m-YSR����( .�~u�����]�ZnJ��J�hM{�>��+]8�>�t��E�����z�����w������T*�Y�������aq�ւrڶl_���F�~�v�ca��7��7�24+��kU.��6AD�(o�[���Em.�d��y�0���0�UV��x�O�Ď���>a�wx��� �J����mE�&��#--d�P��v�,�yPؾؐ��>����o=��#�T��y-��b��t5� ��s�O�C�H'_�s��;��&�f7�u��ޱ���/f��7��M��]��WB�=+Ŧ��$�v��*:��.�d��a���ڴ���\�xobJ�+�[��o�b��8 �������X)�	1w�麫�Ek�vQ����n[M���Ak�C��X��z�9����~�z��v͐ܞ2�w��!�n�:��j�ЉA���%s�?�f��9�j[�	Ź2g��� �����!��ޮR������<��ף�+{)4��q�v�As�� Qh+��8w�0��j�/���+s0���HC&��V�m��>E�j~9Uj��-1|���T�0����d4Bi�i��pN��Q%V��'�L:���"q$ѻ�t�k����z����W�� �Y�p}��p�E����dD��Ү���P�|M�b�P}�y�#
��}s�3u�;���3�k\7��U8Jdz���X���)�|� K8�<`�<��g�3Elǭ���>Տ��nc�oj$��O�=�Řx��������;�f��I�U� t�N�T�B{� ��HD�#kU�&,S���|d :�O�@�޵�@e=��k�n5�Ta/o�#�S�L3ZFQw�����7]g��Gwg6N"2� 8����|G���MO@�����8Lʣ:_�.���=�J�/8wT��ů"|߳�-Xb���݂��OW�2@3/��uHf�U���QZ{W�w6Ϻݔ�5�=kp���qJ>>nw�{F<O�į���[�?��xX��3�vG��ȷgn�M�.�e�vC�_��Q�5?����������ƴ'�����2�D;��8YHڶ%�Ԡ\�n�Xl�����b�V.�X�c��݊�+|���P�.cK�D���Yt�ΦZ�Iv��hc��Qe�E8te�Q�+��r^�V�5 Y�˸�}�_-��b�|���(���`
i*��X�mmc�d�M��
�:����ovJ�j�m4��<��(e-?�yA	�R�+���4�x�;�u��d/'B,TH�bmbc"DJi��Gs�gWq�0�6x7���4[֔�m���)كԾ��d��K����
.�ԓޒQ��R����Y���b^�7�K@���M$j��U,�2�s���	�[���J���*����\��(V��	�s���xL��l��e�uL���`&��p��I��m$��d��j�-	oPz#%G�<rM����-�߃�z�#PHg�O�l1���|����[��)��֋8\�6B}�*F��P�۞})��s�A��!���5 ���n�A�)��[Q��wd�ἄ��3�K����_�� ���v�)����:\\7�6��;���
�^PJz���Ǭ;h��G�s���ᛁ�l\��+��&���>�prv�g4O,B�j���HrI��;�-+x�$e���ja���Dӗk���ϥ#s݄�Z���c�H��7��xK�Ƣ�`�s<Q
�Lbt[����Gd�B�z�~ؙN��O�F��_Q�~sҗ Lb���K������g� 6�:�5���f��M��U{�n�lQ�{w�1�Ԏ�������:ğ������lN��V���~Jq�yk�gx�34� 5��k�֬٪|LF$�p:�����`D��8l��p��Vo
/�*%-�ī�$h�"֌L��̾�(<����HϢ�t�0�Q���d����u0N�ьA,�g�y�Qbj�M����6Ћ�(�M�d�Ŷ�?<3'���k�r�0� m���ԓ��xk�l�n�����,�\���Q�TԴbj��mB�֡$��"���y��@؇\�ܼ������]�:ǟ�~�W�5�zW����0Z 㰧�y�S��j(�8��+Q����a�1�oٳI����3L��� CГ�x�����" ��$7o9VگEA�SN�Q���6O`A�����@6���'��+õ��!�t�f,�_ջ&v�6�*��C,� i+�Ek��%9��ݍC�Dþٸ� ���9~�Xu���Z�ߘ��L��?c� �����㍬� o���;���}V���Et�,Q>���!5
�g����`>I�ӵ�8q�N9q��
�#P�W�U)5�
1�!<T��F�_wVQ�@c���/@�U�= ����~��wV ���w��v� L�3���dQ9#����Ԧe*(E���)8�r;���t��ҧ*O����@���S'󡖂Ҧ����J<�J�Bzw����,��2{���^F�N$RԜ&��ur�FcbΩ�<��Zn~!R��=�T�ˏ^��L?$����qMOY�'Dw��m��]h*�ԜE�t�k4�n�:�6-R�����'rn�{��v��a�9���,����M�`�G9A�{N%�SΩa��?� ����d�V�L1*����b�>�`�I�mx0�i��&8r�{6%���p
�x�I~ � E�����E7[��O��T���l�و�I2�Q�a���V��k���}ģ��>/�Tm�`m.�����u��
���z��y�t��`��G�%Q3z���'P���r���Mr� ���U���<��<�Vxx�Y�(A��t�a�FW#��h�)%8�2o�q�IWL�$ka�Ώ���|�z3ƞE����
o��
Z�}�4>�����6s�	/9��5��%xr쀒��Z��&�����3d�ʹ�Ɍ�Hx串�=�t�6��P��w�����~>��o����MU�9m����� +CKR�Mk.�%)Qpc�Hy��זwD�a�,L��G4:_��=�'ש�m�@ �T��_���ڒ�p�c�F��WϨ ��Ė\�JĘ���{��y\�	RU��h����/%<����������1F@+87
�^#��T��XbF��Ɨe���1��uwp�����|��K{{_��Xl��;P���|�t�UT��Q8�i!��f�Xxi��w� i~-y�e��آf�ju�9e��U�hp�6ṥ4�T~3����]��n}�O�*�J��♎8H�(�c����iB�@`� -��AK
 ��@�� W�&�b��B�H���/�ݿ��v���;�XK��lp�ť�m�s=䘩%�WE7筈3�����=B���x>��x|�9��:Ӊ�j[�{o��l_��Eh�y����͹�(�����"�*d��_�}OD딿�v��t%b��֞�s�ԓ��B�MR���<Xv�x}���s�A��>L�(�U%��I�nK�U.-w^G�|m�r;�R^q��"�kq��J�����"U%65����hXq*{��1�>#d�Gٷ��cfx��z������x'�����FN{�ƛ9������&ձk���fH��P?`��|�3,�2#jA����ywF&�9��^cM9o�c��v��94m;qu�to�?�p��&o杽�������9�-B8�G�� ��.W��\�������E1���4.��Ί�oŷ�T3�����Q�� l���Kk���`�g�Ԇn���O��.]�9h�OBǮ����[O���R��,׹:�/�P�(Q�fY��[��/'���%��G{;.���*�|yߊj��E��P�$d�+%���.���)�L.�@_]�\7�"��9~禭G�1�Q�W/i�+4���Y\��MxF�^��V�]�$.9vnp��C��!`�qN�^}`z�Aɦ<��ݼ�&h��P��>��������y���v+��.r'���RX��US^��5�Q�v�F�4JkE�Tւ�TSk�u��l�g Hݜ����Șm�ǋ��Y l(��)nA���E��h!PGĮ��|�O����]6B�F���,>b |2��
�g�7�4��15F�pR�{ Gk�L.B'4�j��W3J�ͬLs� �yH޲w�=U��N��<]*zc��g�6L5�+����<��3��Wh�%a�) ��=D��ݮ�����P��:�G�&��'�W˽��/Ou��6h}I���X0c��������v@v]��.�X�'���K,�����;&#���w[@�L�0�r}���j�%���5�L�P�(�(y��U�E;�T�A�~���c3�����$˫o������e�4Q= �����V�GUZB����ӳ-�B�����SM5����I TKC�qN*;+�$�˝~�mE��yȶ^�K�V��q�u{�XT�>j�<do�u��-YXi�*#����!>�6,�w�B�����%�������
7v����f� ~�氷t���-�q��nw�]�HN���mo@|�C���|}۹����A����6�$�/лmK.��8ھ�V���~�(��_4��E�ֈ<I*���H+��ރ���������ْc�fPPOn�#cID�����E�)X](bȺ%6(%nŻ�́�\sk|��
��?�Ò�0%���֥A�HCau�٠���籇P����.O����k�?_�K�5��F��U�'r���ˡw�V&���S��Ll��L����s�B2�.tf���I�닎��5�֓z������T�l�-�B,7�A���a�a�����.H͛�xcn5����F�F~9�����ɶl��]���hj*-3@t����<�7�7���[л�w/ui�fj�/�|"!��y�MaJ]�Z�ᳪ.e���C�X����*ˋ���SI
��H�
:�v&aEHA(�Z�ڒ�sR�@��..F��H{/�Y
��ڇ�Qad�q�0k�)���>��A(v.h�I&#���W��q_dy��[�������ʛ�ͣ��澶r��)�*T��u�T�+1��^��2�<�A���	��t�oי�N��� �W �ˌITv�J~t�)a$1fw=PY�~�d=V׋��ea�>�#����
��"ə�`�G��,;+C���_��86��ܓ��L�� Kz����J��a�+�{�;I�w��=a����K�����dG
�Ibg�Xl��ݠ���m�ʈ���mʳ�3�Ȏpn���`nJpS�&�A�����&=)���q鋨��e�n��8�e#@.���u���}L3���HG� ���P�a�>�4p���\p�S��J�YQ�c�W2��,9�g�ז�~���I=tx�¢߲�m��4�f��\.U���� ��esQti��Z��5+R�`ĭ��YD���W1�_0�����(ЪK��Z��C�"2 P�V?�����#4+�o4c<���D�}�O�m(�@X�~��,[�q�h��J�d\/Q��GWE���L��V�rG̮�4svL{蜍g.���\��g�^)tĜgW�q�|�L�.&C��0��/`΢�lэ�-Jb��R���a-�_��I�X��j��Ji�&agy?�)>-�5A��Bc�W%c�h/�];WF�7�N\�=�Q�-��̮��s��4o���(+�
�4����4�v壂^ņ��NH;�3����	s��ݨ��8��ɒ_g�����!2����AqF���R�` ("4�	8oK�}��68\��i�lIQQ��g��İ��+�j>o��;U�m��/^F�a#jl��,gń�H4iUL���!��z�Y�ڀ�ׅo��R����J,��$^�z�ɋ�uy$Q�4���b��z@��� u�z/�I�����a!tY�vB�On9�m��/���� �5����8���iF�zY��ǓЧ�͖��Jmq���YI�z�R�l@��g��N����0j3{]��2J[�ی�
�Du)����B��	�3�Y���%�29�o�q��N��N(��F��}L����^2����5{ܪ��-2���y\-��?w�����C�X�׫L���+�d������]��P�kl*�gju'P�Ea�/���	�r������ّG<6�#��k�KW��R
0jG���v� U�+Z��
q�8j�����4�XO[�5��.�	s��������h+[�#"�����7f�����{��<�)��W+^�#�5�_GwYl������){����7mÜ�D�ִ���ԱX�;П���J$�7��[C-x�
����s��&���!?�1�	1��)e��"*�81��?ZX���F0h��<��P��2��H2Xb��3H��[���n�(~��f���R��0'�J�5<�6PvY�U�{j�����]�Ȣ��
Ȥ<�r�����������<���X�xۈ|	(I���F��9[���w�0�r�ʕ[i��V[�si�Qh1�a�/1�_t���?��~-��T���EsU��FY��$�D(hD�R5�?�		:�K�`��Opq��w-�k k���?<���6\��u����x-�~xb��5�*64��ю�%Ӷ�;��t�K��_�ޓ�f�9���v�`M��~/��aV�y��mG�E����ͨ�@�e�6h��8�o��=$�Ӭr��T��i����O��)�m ��b��U��*�=�9oj�8Ō��8�β�GbLb��}���\���t��t�����2��ΠU�o��OgV��?������Fxn]O,c���^�~_��aIFLi�.nQ��O㯐иT|W�I�O}�^�"=���*��a�l����ﵪ�Z9�P� �[�AzM�ҧ�b<7vE�/�k�}�nԻgD}������^���p�M^��QQoO�G��.$?�4�ň��䜍��l-H!o��^/��~'�)�ԇ��������e�w�v����PL�7����?%��k��ȣS��d������"b��o��bձ0�zs$S<���
���I�b��[~���_.Wt�:d[o��qԺ/����+��ۆ��[��?g������^�H��S�iw�"c?ZI�U�-Ȁ�Ų���*���hi�`��A�
&�`3�Yծ\谴�,�U�����Ƚ��Z���� /���3�4q��=V�	��qj8�OS�_��ξ��`F��`������#�f:V�z^����}jy��9
c��OnB�`t� ���l�gK����sXָ�y���A2χ(�V�FhԂr�0�}<�>BN�8[G6���[B�<e�Vmz��5M��ꐜ˱������I�ނ��OR�~�r�P�
iZ$�i�Ҽf��RԲ'I���^�0TW� 4��XY/-!,�N[N~S�Gi��'Յ/��f��ޡŜ��I+����g��4�@Q��?��(���~�C��V���6��jfgS������X5O����R��}��M�!�Y��R���Ep����>�WBwX����>�(,e��X�в(�/2#��+R)6W%�Ĉ�Õg8�|�B������
�"�\�����$wY�y�)���ANմ�wM^B���#��qgk��"�b���=�ɷ=쏜EW! �4����_�����Z���*h
s�5���d
�Տ�����k��R��쥙��Ϝm���l��^zx�C����ز���]�&+/f]ex���j?\�TD��Ԝդ}O�ɕ^h YP�d������L^�t��ڭ����GON�8�5�Cŗ������`W��^4�B3߁v^��~g2���Ő�F�BR'�K
�.�+P��k��<���/�y��E�Tu'�s_���H��W��=f4s$/�^���Q`Qe�}?���l�B{����h�#_آ1.���{�n����Iv5C���%H( �b�%�  Ӊ�e�r��76���8����K�/�6 �Q0�f���i�g;#
W:s���b]B=���p�����MmJ�eiL�k��6�5�
��4C�}�k}V�.!GZ��H��rqܝ5�����Wk޼,�	�+������!��g&i�Ƚ�B������Ω�a�{wY��w��KkL�>�%:A�8�)�bJ2/���Sa9soyy�$'���
+T4�Yn�$gf7�D���W��?o���<������bO���&�S�GJ������A�s�__A;�i����^��4���ԅ9��FL�U�*���?�?� a�1hI�Y�VQ�Di�#ZR�hi8�����c:����U����ڣ:�K?�z"�q6��ₛ:����wÆ��q�Jc���z�ߩs���������b��&��[��"����V4��T|�u8�1�<y"g��I�Y���T��c������Bd��r�}�%,�?%��^0սyk��x�:'��v��J<.)�Ԇ�R�����IcD�ߕ^g��&�b�y��?[G  �5OZ��X���d�.�)tIwӵ�yێ��ݩ�����u[���(C5�7��d�-4`�3j��M*�� r��4x�RI�>�n�xp T�a��Yy��Y�^7"�b�[9���Ar�RKR�_�>�v<��g���K�_i\S��RK�PS���_�g��
� �Lh���(�&$���CpN ���1n"!B���^�]�l�(�