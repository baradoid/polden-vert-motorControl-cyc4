��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�=l��!ӻM�׬�d�#�z�%8/�=s�oU`�&���g�$�m��^����>���ŉ����;��= [g\���{ b*Y�����?mX�L%I�uG��hB��>�ED-9�8�����6c�>����쩶�X�I;����]S��GP(1�OAk�T��{K�9QO�K�����S@o3�'�%r2e2W�${满!��b (�$0��������|8���+5�p��y�F[H�[����.�1Ռ+�~�����s �Zɷ��SKKZ|�����`�|\��`\�!��|'�ö�WOY<�$�8��N�BF�F�B_��f�a[�3�����v�X[����l#������N�-�A��3E~�Ye��&Yʭ#�ד����[�����������@B���h�i���Zk�-���<�Z�M^��b�d�s�75��5�	���3���H_`�A�E&m�5I���C��ܷS��T�������5������kQ���T˯5=ԅ��j��[��M���0s�ud�~z���l�BOr�*�/ݧ���,r���Zv="w��D����+;4o��S>WE�>�k�K��I�Q�c�p��Qx�_����!Ǌ�D�-�䖠C�>��_K�7 ?5��͇*#�IY��h�|��»��y��y���xc3�#)n����Ux�M[$eh್f'�慕��kj