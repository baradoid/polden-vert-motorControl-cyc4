��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��[���^���3����UA�p]kB뷜���lo��2��6�5�F�=����D�:jz#���L��s��u����}�9v��Iያ(��p����ðT�)�O
���� Q�b�&'�4e�x-s&:�V��c2�uo.� �o�{�r9t�����mZs����SҟN.q�֨�&OJqC{�.�ԍ����I+�4XD��P�,���p�AD,��[�]�*# ��HI$ps�{^=�����A�6�H
0\���W���䕮�0�ȶ�@���E��m;�в�l
9
N�l��9�0�D�uR�T��Z���h>�0@��A���QWg<����y���!�g8��E�������T�lM5��@¡d|�h[ȋ�^��y; 2z�&�����ˊ���xB����U=�0��ɼ^/��L��t��kOR���C����xF'ZN<�Da�8�\r�Ri
�(0�`�C�2��v;]�x9Ukv��.zb�;����>Yd&9���C����������q�l��*j�2�Ҹ�0%��D�`g-.���v8�����������#,�2�:h�����$�G��Գr���c�����?���y6�w3��i��'�K)�M��6^i��d��E^f�T�~��P}��tX<[��[�GĀ�<`�Npc�ɸӂ�o�s�M��e���uJ5���p݋wkY�B<�]�x���sOyq6`���ʴ�&���V�������3K�v���d(���>�"���I�~�����cN������"�\��o�I���E=>c��g������g��$ �$`�t�va��27Gsh�����?z�u���j��ҧI�J�zEg����e~��`E���vsV�̖t�˅�dYR�+����Pd49����q���h$e���0�L����:@���*��q�RehK��Ƌ��zM��>[ .K�#.f?�6�ks��-o��]��,c�G׵�绂�Z��3U���λ%
��X�347���S�禺QѦ����-��8o;�U�Z�b�m�	@���(��ޔ�ߚ��" ����y�O���G�.��h���6��k�c^l�c�S{bS
�U�n��vL?Y��
N��Fl{B�?��ofҿ��=��4�v�ҹ�bT�$a�d��]����Y�T?����*�7Ď5��<7Mp�[|>N�$���M�,%�Cs�{����i�r�ɔ��J��o��&��@�F6�u6�)$D=��q�U �k�������+a_���<[�����}6
3{c�pXl՛&�	
l�I��ؕ��F�\4qx�� �Y�����Љ�0�h��F�r.�MA �	��i����KbU��:�{D9x�5-�0�J��2���	�F����Y5/OM�P�|��Xs�eq��Qc1����p`������.�S{Rj�bهR�;�y�h���͑�Hg�%��P�g�u��JD��
I����2��Y7�.�#3\��#������]i5���4�;[pQ�#@��>*C�ȥ�L�^^B"�F���TT(L�#��5�X�����J?2L5���w��T� !Q���JN�"J�A$$��^�2�^�ʂb.KO>����($��6��5��2�dJZ�.^�kQ�e���4g%8���R&l�Z5����} $�:(r���z@+�m��E�inWQ���|�S��c�$�E����k^ @8-��Z���K<�ȿ��f�[R1lѝ-��U◖��gM�����z��2���X~��4��u���&�̒�R�蕯x�P����d��﹋S\�j�J|�ªn�S���r�@]ul�e&VH�v<ȿq�6�Ʒ݅���]��0�E�L���K����a�îY��Ģ���6|c*X6)���*����+�zl�q텫P�����d�˾]h����n�~H�@�r
��мEX�`�ȼ�<0�X8�v��K���dԒo�͓�L���'T䨝~(�%':�^�אR�k�K|C���m��ݾm~�$�O~vM��h��������*G��|�iG�|�$]Nj���#�n�!?���.�I����=���lF��BFֈ��٣��5:�W��#���
����5C�2Ǯ(a��:����K��C3u��v��\�'.�4���X�2���� �Q�e#�I��g^���^k��T��Y�=�K,����a�Hʍ�n�m̕��,�<Ы�=��`�+��q��]ǭ�;�%a �	+؆z�S.�w�1B��� �Rj�GS�L)IeҖ�U<���ls@t���'TɪXI��^ɰo��K4_�-v���d��{�����z���M���4��6�ʸ�d82~F��+<°��y�
	�ɂ�.$8v�)pY����VI!L?��d)�ֳ��l���H3��mx�U�Hu	�Bo@��/Hl�m�G���%���,]�={�Jpxab9]���
J��0��`o�a�}���[@��!�PUa��c`*Us�gX�յaT"�o����l��&G�]��2�;@4"m�o�1X��?v��C�B/�^���.���[��U.f	eg��g���h)(�;�VrHn�)�(��G?w�V&�3K�eD��Q)�i@?�f��i�DktI�tѯɗĂB^�ơ�