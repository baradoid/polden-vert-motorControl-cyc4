��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��[��F[����w�g�	�ɞ�/8�~JE��ƣR��,�gU�j���}�~�(ͤ�5����[�d��r���v�W>�{�~�@'�G�[����;0cV��:������An���?{#�
3���������EA��G��,5X�� ��t0HÆ��]\�DX��o!��`&���/�3����/d�Sf	��1!L���i�M���5��p��Mw�H"��!�mj}X��R���*���:��Og�R#���-�����KƱ�q?Io��D>՞���p�'
bIŰl�jK<ϔ��D�l���#�)�V.R��[���ٝdJ��6縪)3��1vt9���$"J;���.��A�F�°&\�?r˫�;�}�?4j]rޯ��/�C�"oK������Y&�_:���x<f�,*���n���>�B�i��s�pax��=W��A��+�K�\yq���#"�����t��Z!�s-�	-?*ƣ���'H�7�Fq����S�1��￐*u�ʊ�Ǜym��O�Ģm�#��}j��>�dK�����!���X�Gw�뿝��Ҝ^yV�$���١v<ëŭ��q19���.���r���.��0� /<��7��Ӌ��2NN�X+��L~�Թ��Ы�����MNu�qQ7�G�A߯�{�#^�������1qצ�H��=����]:k'�+jTED�Z�e6���b�@|,_OF����X�������>T`@�Ԑlw�1a0��Ĥ����5Zsκv�S���MQ���(;�;�oT\�Bpg�Uˊ���0 ��8-Q�o��܄p�3{�@��SW�ݯ�11���tD�{�e�$b�6d�=�# ��k�A����P�	Ϋ�g�v�­l�b�t����c��[�l������V��M�ξ3���4Z 0�ިʪ�Z߼K-.���t�r'G�~Ԗ��\e��6L�X�S�b��EI/PQ�����Y�
��1VT@N&yy��z��X!y���W�Þ��(�(�MHD����훐�#�^v�T�/'�Y�v A���~^��	ӽ�{lB���e���	�$�b[`���Il�k��a����<�H�vϖ��l|�ǅ�V��!�H�[R� \m��
��T���%��3�a�P�@L;,�����謌q+ȭe6���"p�HT�Q�C��X`(@�Gszsh���lh��@!�kv���m&T{[!K����9Z�qP��c�!�˂��d:�'y���W���;
�J�(�Ȝ{��UQ�dN����Y|fn�|�>���E:*<�N!�[0�n�_�ӽ����	K��&|WAZ9���'S^����ɲsx�5=%hT��#��c��C�S|���:�.8�����<$��-�ޭh<��'������P.������ir_tE6(�|z������D�ج/Z�/��I�0�X�<0�@���/�88��Y��`P��5�d�mX!�0	>$C���kN姍��ߑ��jۈ� �y��Y�ٛo��ǽ��邏E>6Xa�$^|MeVB�BSwVrl�A�������A���0�R��_`�w��߰��Tr�.P����k�{�&)~������*_�ς���B����T Q���z���؋��'�h��B"5��ԏf�#�a�?�D]e਒���h
e��m�DD�W.����/U����t31�j}�)� SYuC�k ��"=7�Yd�S�3��=q NJ��mq|�Z��P��x����7��i��C�<�侎�c�q�8�wE6֟0���w/ ȵ���IP0����/��6/�8�>� ����0E���~?�m��
�Q�}箖1phShx���f� ����/)I��G�2��{�(�-��ɽ�����◑NI%�}%VyI����A�!?�@��IԬ�V�m�U� C &-��9���[�/2ydK^��(�V�u�r�0�%���TwI��V��:�SX���B�.説���ڴ��g���-G��,~���i"G��'T厩�%�	���7�V��!�x���ٚLi�w)��G�2�>�]�H���!��{���p'�V9�Փ�͠����S��Qr��`50���6�1�b�G�:��	2��H����b@�VD}�{r��{���G���ú�1�k0�G`����B`kZh�F���l()׏Z���/N�%�>��E��s�gj��6B��7��Ƣ��kYW�F�u:�}g_�E!&F�J"J�-�C�7�ߩ�����Ӈٮ��/���3��#A3�uc���eV�Pj���> �n^��5���tJ	���.�@EUA�(jq)�m1�l*��a�Is�onr�I��;IX�5�5w���͆�	�P�6�ˀ��B���P�MK�~P���I��T~v�d�"�� k�o���f�X��)�>w��G�`��tv/�w�c�i��T�~?9φ����7�g@�[�[>Y����p�Q-������)��h���x�p�"V�X�o�0
��=��pdɨ"��Y �7	�	f� }vV\g�M�A���]J_���A#�K0�IlO"G/2�������ٷ�m��3{�|ߟ�ك��oi�*3D"�
Q�\h7U����	����w��������M��6^5��� P��21���P�֧G=���z�8p�
D�c���
���j��a+3����p4��r�D�V� B���8j�Μ�i���`h��pU�cg�Y��5���?l���G6ԅr :��d��(s�I�['��~P��֨m��9e�@D�6m:����|���S�!%�:��[�1��*��ߡ��a�A^gWql�9�<U�f0����|�5�5�{}�6��C{�0�D���C�VA��|���q���r�p��g���2G:�x���K�������^�\G�����8��� ��WN�7���EeM�|[T+����e���]K������6FEgn�9�@����}ʋ�B����_�s��_�A.���&��lU׬�����Y�>�4v �����r��x���axR]�'U��S0Iz���a	,@��*q�Ha8�i�_hÛ��E��6��r @�v���sD�k����4��qH_��J4�%v�U�'<���*0m.⮦�dX�c��yV�"J��S]���)d����sA̺I�D�[,?��ut�uicG͹�/�E�(��
AcF��ީ�Bɡ�R��
2e���m�Q�3��N�A+%���1�ho�ܞ2�MO>3n�עԄoE�r�c#k�m�(S�7��C�O����j���T
��cax8���/|<�#<{:��N�"e�ݾv�����V,8�����inS��=̨�2q�ٟ���+eϕ|�U�Z�ifiZ�ā��F�@�̡��e���§)�!��A��"wU�Z�"9�Ke��.��q�!9���~<��^��8�\����`{D�� ���c�	����"bu�Sr=��C���QG-]O:@I������yl������;Av�g5�K�\Z���NWf�ч�ڴQ�_#x��dC`UM�T[�y���cF��^�Ai����5��\�'&�Ǣkl�