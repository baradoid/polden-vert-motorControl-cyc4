��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�
#��.{иp1��j���HX�_�Lqr�����}�Sw��n5��p�{dB���5� {�@��b�·�I�����:�S����UeRQ�c���¥;� a#t]�?����OR\��iY��Z���]�߬�F"���K��j���႐$��f|"��F�H�_� �����(k���+�\��;�|v�E�+xCڬ������GS�p��*���K/�3�]�M�$�7�k�"Û.	�'M�ƹ�u��)������%�{��&s7���4\�����*?�I�!��z�47�V�/�sO6���,BTm�f@��4J��F������|qR�qZɧz�F͎�A�fQ۲/N16X����K-�t�&1ז��6�(݆��X_��o�&������KR�-κ��Q�<w4ڀr���\���Bh�q68��N�ZW�@��t�kO�Tc̢��K6X��z���,`�f/^�_)[�~ ��G� ͞h��e&���-���e��ښ��Kɻo��F�M2Zv�%�3P���y;��ng=)}*eDu.f����U�˸�[���Mmd�C��������}P���+8�_�[����y��hx_����o�P�q4��'U�N���������=Ů��gf�$����<���V��DH:;�-��ha����/�!�t	�n(`&1l���y���v'n���4����������Q~����v_�Ӭ�,��Yxzun~���G��Kª���7M�K����ß����1���~91�;��;�f���&�D)���_���#E�����_�����P�s%��}�A��y�zǂ�0䧒 Xg6��6��o���[2��+�r���wB�V!�tz��s�ˎx5�ij:�J
����?��u>Zx�=���&#�g�Rˊ5q�/���v-��l�|�+oN��� �xk�iPO_�Mt��LQ���w�hd���b#�$ؖ�C�AX��F��O�F/$I��t0�곀���+
QW��쬵��ϣ�����iBL�}��������q�g�s��[4��L�/��n���ΖZV��'_\�:V�l]?�2PH4�E��K��ءhE��'�ƍ�.��y1�-�
����o��D�V�F#L�+ A�бG^O�'����pz:��~��*n�ػ�>Rea�㬯&T궬�D��t��ŕ�A��"��a�Xd�R����� e���za?�����O���o��~\[��MD������YqI���P`G����E  ���T�&�hW�k;���b�4�� �A�e�O��U �<�m�`1ZI�>2�c2�$���1��<�Iȹ҈!N
�xU�{����i��#�R3������S��F���؍��b�e��G��Y�ҿ�n��Y��SK{��Ix�(D����c��o5�$u+a"~�?Wx&��Q3MWu��܃�����Q�|���/������������\�.=�f�B��y"9�Ή����<ứ͔4��BpB�\���oJzř�9ˋ<��v}"Ʌ��.>����´	\-���l�.Ǻ��k�n�G��~�T���|o��N�!��8��ȁ�zE��C���w�4�E(�6x~ u�h8}E���e�"`}�p��cI���q�ɸ�A;0���#$:���������$�]w^dϝ�S��L#*MT��<!(�!�N�����z��Ǚ4!�[��Õ���ޝS�|�9v���?$��Ԅ�Dg.&+��wR)w�;ɵ0�]oJ�,'�YTmYQ��-Q�:`�[��3�͏ ��V 9�w��&6$g���r�.��$���M&Ɏ�TBVꬤ�=�/QoT�ʥ{�+7ы�@�,�3�7S��8!��u����}���k��r��
��e���K%�Mג7LM��񯡠�l��l,<�L�j��c4���s��֞.A�{�p�_����@�eB�&�:�)D�C�Dw@4@;O�N����Y��B��G=;�CxK���9�<�v�4�<q�}���E1��3�b֨ox�_E�$)�*��x��Z7���A�Z�a�	F��Бs��.����"S{�������	G�9��D?ΰ]��##5���>fl����y�%Ai�%e�%�E�G�(��K��M+�Q$���W�� W�}<B���R��y���e,�l��^U�6�Q4�J�5��2��t��$�q�Vw�ץ>Ȧ��%�851�ܡ���m�2X*�*ߓ5�Ğp��T���z��Y��^��=E�,��n[*%bm����TI����W����j��jݜ�vc>���ӿ�y)��$�ٱV�"�]�[A�ݤ��6	��CB�nc����i������o�h@�K/���K�R�Q������
�������|�g�/+2�"��XF������^^��ʖ$�U�x��ۃ汼9\*J��UXOg�sB�{i���������sC�ݏ��=�˸E��'\ސ�텁A�{O?~q�G�6�NZ@;V��`��bJ���B�����w�pP��L-�G����@�q���s��]g��o!�����{>�>�#�Z�f�[�Um��
��q���=�OY�i���	ZSl;��"�;� ���u����9l��.��n��ᯋ�����گT�k�H ��H@��eD����I�[_J�ck�<n!�EINJ�:-Q��[�,���ڕ-�(:��㔵�?y([p���Vb�ɥީc��b_Xb�I�<�����~J��z*��S�^sD'��%������0Q���Sh܋��Jޘ=���=u������U�,��z+����~�!x:��s"���D+��wY)���q���^i���q4���a�c'�};�A����u;����H�o�F^D<�fE��N�����.{Ce������<����`x��j���e��dT�9�A�����ꐚz��w<��d�od(S%L�Îԍ�֏�uI=�-�㑷k�KMƋ���$Q4=GG���ۉ�煹f!���?�UHq�l�^����9���q�[=�3����r�"������	�ȋ���Ct��-{�S�;`����<6�Q~��У�y�@�>�����;�rRŽj������Y�ss��d�O�b�2��z�@���k�m�K���o�S�ld���k^��.T1��w����������ZZ�����U�����W��:M3a ����#���r��Y\�����V"$׆(Pλ��@�:����ϣ4��S��HZZ:������v[�����GO�|��U��f����
�����Ζ!/`ƀ���R�����Z��_�)0�W��k����M��ZI��:/�%z�Пr��+��fT�$qɘ�6%�i��؁�{���c-
z�-��⾰K�&B����>��_�3|�T�������-��{��J�XS�^�E��`�J�&�Skcn��:EM�-AN�y�#̿`�r�)\����T�<r����r��Q0e{��v5:ަ�@f����S���e?i^T�!!�Q�"�;lh�pÓ(`����&��؝rb=�������]�;�lRd-Om���9��#P�����	���r�Y�n^�)j���m�
'B����̵���Nt:X�E�;�`�⅕x�����s��QWS�<�"O�ہ.�06zܟ���挒s`��{.��fS<��ް�f�t���[��n��7=bv�S�%>'#8/����Y�)r�}D��!�Κ��\8�w��\'"H�R��	vQ(�H�,�o��SO��2��΍Tk5^֕׃>[�������$���b5o�8��c��k� I�a-�k�YY�-���ݭu6�ֽ�AQY���&[�=Å�dL��l=��:LdUG�6;E��M=��¸�7:�aō`�#F�yp�,�/D���'��)�@�.�E%�iV���m�*| �gٳ�`�n�6�"tB�w�<�Y�3�rK܎���4t��ޔpjb-cmL�֑\�� �Pٔ_իEGٳ:![m��7��7�z�6�)�O=X#CՆ�CC�Z�Ρ�b�Z������������ŴOX���q�R+���E�+����R���|#������C>��a߹�p��)1	�i똱{�ׄ�[�~�
�i8��zG�